module router_type_2_netlist;

endmodule