module router_type_6_netlist;

endmodule