module router_type_3_netlist;

endmodule