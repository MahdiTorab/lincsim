`timescale 1ns/10ps
module sv_router(data_out_array,
                 sent_req_out_array,
                 new_out_array,
                 ready_in_array,
                 vc_no_out_array,
                 data_in_array,
                 sent_req_in_array,
                 new_in_array,
                 ready_out_array,
                 vc_no_in_array,
                 busy,
                 my_addr,
                 pe_id,
                 active,
                 reset,
                 clk);
                 
parameter each_cluster_dimension=2;
parameter cluster_topology=0; //0:Mesh, 1:Torus
parameter cluster_first_dimension_up_bound=8;
parameter cluster_second_dimension_up_bound=8;
parameter cluster_third_dimension_up_bound=5;
parameter no_clusters=5;
parameter cluster_first_dimension_no_addr_bits=1;
parameter cluster_second_dimension_no_addr_bits=1;
parameter cluster_third_dimension_no_addr_bits=1;
parameter no_cluster_no_addr_bits=1;
parameter have_fork_port=0;
parameter have_express_port=0;
parameter no_outport=3;
parameter floorplusone_log2_no_outport=2;
parameter no_inport=6;
parameter floorplusone_log2_no_inport=3;
parameter no_vc=13;
parameter floorplusone_log2_no_vc=4;
parameter flit_size=1;                //In number of phits
parameter floorplusone_log2_flit_size=1;
parameter phit_size=16;               //In number of bits
parameter buf_size=4;                 //In number of flits
parameter floorplusone_log2_buf_size=3;
parameter switching_method=1;         //1 to Store&forward, 2 to VCT, 3 to Wormhole switching
parameter addr_length=10;             //In number of bits
parameter addr_place_in_header=0;     //bit number in header that address start
parameter [3:0] my_type=1;
parameter [31:0] node_links_directions=0;
parameter want_vcd_files=1;           //0: no vcd file generation, 1: vcd file generation
parameter want_routers_power_estimation= 1;   //0: If you don't want to run Design Compiler flow to estimate routers power, 1:If you want routers power estimation (guide for more details)
parameter is_netlist_provided= 1;             //0: If you want estimate routers power and provide netlists set it to 1, else 0 (guide for more details)
             
output [(phit_size-1):0] data_out_array [(no_outport-1):0];
output [(no_outport-1):0] sent_req_out_array;
output [(no_outport-1):0] new_out_array;
input [(no_outport-1):0] ready_in_array;
output [(floorplusone_log2_no_vc-1):0] vc_no_out_array [(no_outport-1):0];

input [(phit_size-1):0] data_in_array [(no_inport-1):0];
input [(no_inport-1):0] sent_req_in_array;
input [(no_inport-1):0] new_in_array;
output [(no_inport-1):0] ready_out_array;
input [(floorplusone_log2_no_vc-1):0] vc_no_in_array [(no_inport-1):0];

output busy;
input [(addr_length-1):0] my_addr;
input integer pe_id;
input active,reset,clk;

wire [(no_outport*phit_size)-1:0] outdata_vec;
wire [(no_outport-1):0] outsent_req_vec,outnew_vec;
wire [(no_outport-1):0] inready_vec;
wire [(no_outport*floorplusone_log2_no_vc)-1:0] outvc_no_vec;
wire [(no_inport*phit_size)-1:0] indata_vec;
wire [(no_inport-1):0] insent_req_vec,innew_vec;
wire [(no_inport-1):0] outready_vec;
wire [(no_inport*floorplusone_log2_no_vc)-1:0] invc_no_vec;

genvar i;

generate for(i=0;i<no_outport;i++) begin: outport_loop
  assign data_out_array[i]=outdata_vec[((i+1)*phit_size)-1:(i*phit_size)],
         sent_req_out_array[i]=outsent_req_vec[i],
         new_out_array[i]=outnew_vec[i],
         inready_vec[i]=ready_in_array[i],
         vc_no_out_array[i]=outvc_no_vec[((i+1)*floorplusone_log2_no_vc)-1:(i*floorplusone_log2_no_vc)];
 end
endgenerate

generate for(i=0;i<no_inport;i++) begin: inport_loop
  assign indata_vec[((i+1)*phit_size)-1:(i*phit_size)]=data_in_array[i],
         insent_req_vec[i]=sent_req_in_array[i],
         innew_vec[i]=new_in_array[i],
         ready_out_array[i]=outready_vec[i],
         invc_no_vec[((i+1)*floorplusone_log2_no_vc)-1:(i*floorplusone_log2_no_vc)]=vc_no_in_array[i];
 end
endgenerate 

 defparam router_cortex.each_cluster_dimension=each_cluster_dimension;
 defparam router_cortex.cluster_topology=cluster_topology;
 defparam router_cortex.cluster_first_dimension_up_bound=cluster_first_dimension_up_bound;
 defparam router_cortex.cluster_second_dimension_up_bound=cluster_second_dimension_up_bound;
 defparam router_cortex.cluster_third_dimension_up_bound=cluster_third_dimension_up_bound;
 defparam router_cortex.no_clusters=no_clusters;
 defparam router_cortex.cluster_first_dimension_no_addr_bits=cluster_first_dimension_no_addr_bits;
 defparam router_cortex.cluster_second_dimension_no_addr_bits=cluster_second_dimension_no_addr_bits;
 defparam router_cortex.cluster_third_dimension_no_addr_bits=cluster_third_dimension_no_addr_bits;
 defparam router_cortex.no_cluster_no_addr_bits=no_cluster_no_addr_bits;       
 defparam router_cortex.no_outport=no_outport;
 defparam router_cortex.floorplusone_log2_no_outport=floorplusone_log2_no_outport;
 defparam router_cortex.no_inport=no_inport;
 defparam router_cortex.floorplusone_log2_no_inport=floorplusone_log2_no_inport;
 defparam router_cortex.no_vc=no_vc;
 defparam router_cortex.floorplusone_log2_no_vc=floorplusone_log2_no_vc;
 defparam router_cortex.flit_size=flit_size;
 defparam router_cortex.floorplusone_log2_flit_size=floorplusone_log2_flit_size;
 defparam router_cortex.phit_size=phit_size;
 defparam router_cortex.buf_size=buf_size;
 defparam router_cortex.floorplusone_log2_buf_size=floorplusone_log2_buf_size;
 defparam router_cortex.switching_method=switching_method;
 defparam router_cortex.addr_length=addr_length;
 defparam router_cortex.addr_place_in_header=addr_place_in_header;
 defparam router_cortex.my_type=my_type;
 defparam router_cortex.want_routers_power_estimation=want_routers_power_estimation;
 defparam router_cortex.is_netlist_provided=is_netlist_provided;
 router_cortex router_cortex(outdata_vec,
                             outsent_req_vec,
                             outnew_vec,
                             inready_vec,
                             outvc_no_vec,
           
                             indata_vec,
                             insent_req_vec,
                             innew_vec,
                             outready_vec,
                             invc_no_vec,
               
                             busy,
                             my_addr,
                             node_links_directions,
                             have_fork_port[0],
                             have_express_port[0],
                             reset,
                             clk);
 
always@(posedge active)
 if(want_vcd_files==1)
 begin
  if(my_type==0 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_0.vcd");
  if(my_type==0 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_1.vcd");
  if(my_type==0 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_2.vcd");
  if(my_type==0 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_3.vcd");
  if(my_type==0 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_4.vcd");
  if(my_type==0 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_5.vcd");
  if(my_type==0 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_6.vcd");
  if(my_type==0 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_7.vcd");
  if(my_type==0 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_8.vcd");
  if(my_type==0 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_9.vcd");
  if(my_type==0 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_10.vcd");
  if(my_type==0 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_11.vcd");
  if(my_type==0 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_12.vcd");
  if(my_type==0 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_13.vcd");
  if(my_type==0 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_14.vcd");
  if(my_type==0 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_15.vcd");
  if(my_type==0 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_16.vcd");
  if(my_type==0 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_17.vcd");
  if(my_type==0 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_18.vcd");
  if(my_type==0 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_19.vcd");
  if(my_type==0 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_20.vcd");
  if(my_type==0 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_21.vcd");
  if(my_type==0 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_22.vcd");
  if(my_type==0 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_23.vcd");
  if(my_type==0 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_24.vcd");
  if(my_type==0 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_25.vcd");
  if(my_type==0 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_26.vcd");
  if(my_type==0 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_27.vcd");
  if(my_type==0 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_28.vcd");
  if(my_type==0 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_29.vcd");
  if(my_type==0 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_30.vcd");
  if(my_type==0 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_31.vcd");
  if(my_type==0 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_32.vcd");
  if(my_type==0 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_33.vcd");
  if(my_type==0 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_34.vcd");
  if(my_type==0 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_35.vcd");
  if(my_type==0 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_36.vcd");
  if(my_type==0 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_37.vcd");
  if(my_type==0 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_38.vcd");
  if(my_type==0 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_39.vcd");
  if(my_type==0 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_40.vcd");
  if(my_type==0 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_41.vcd");
  if(my_type==0 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_42.vcd");
  if(my_type==0 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_43.vcd");
  if(my_type==0 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_44.vcd");
  if(my_type==0 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_45.vcd");
  if(my_type==0 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_46.vcd");
  if(my_type==0 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_47.vcd");
  if(my_type==0 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_48.vcd");
  if(my_type==0 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_49.vcd");
  if(my_type==0 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_50.vcd");
  if(my_type==0 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_51.vcd");
  if(my_type==0 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_52.vcd");
  if(my_type==0 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_53.vcd");
  if(my_type==0 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_54.vcd");
  if(my_type==0 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_55.vcd");
  if(my_type==0 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_56.vcd");
  if(my_type==0 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_57.vcd");
  if(my_type==0 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_58.vcd");
  if(my_type==0 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_59.vcd");
  if(my_type==0 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_60.vcd");
  if(my_type==0 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_61.vcd");
  if(my_type==0 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_62.vcd");
  if(my_type==0 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_63.vcd");
  if(my_type==0 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_64.vcd");
  if(my_type==0 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_65.vcd");
  if(my_type==0 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_66.vcd");
  if(my_type==0 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_67.vcd");
  if(my_type==0 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_68.vcd");
  if(my_type==0 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_69.vcd");
  if(my_type==0 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_70.vcd");
  if(my_type==0 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_71.vcd");
  if(my_type==0 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_72.vcd");
  if(my_type==0 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_73.vcd");
  if(my_type==0 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_74.vcd");
  if(my_type==0 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_75.vcd");
  if(my_type==0 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_76.vcd");
  if(my_type==0 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_77.vcd");
  if(my_type==0 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_78.vcd");
  if(my_type==0 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_79.vcd");
  if(my_type==0 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_80.vcd");
  if(my_type==0 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_81.vcd");
  if(my_type==0 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_82.vcd");
  if(my_type==0 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_83.vcd");
  if(my_type==0 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_84.vcd");
  if(my_type==0 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_85.vcd");
  if(my_type==0 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_86.vcd");
  if(my_type==0 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_87.vcd");
  if(my_type==0 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_88.vcd");
  if(my_type==0 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_89.vcd");
  if(my_type==0 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_90.vcd");
  if(my_type==0 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_91.vcd");
  if(my_type==0 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_92.vcd");
  if(my_type==0 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_93.vcd");
  if(my_type==0 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_94.vcd");
  if(my_type==0 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_95.vcd");
  if(my_type==0 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_96.vcd");
  if(my_type==0 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_97.vcd");
  if(my_type==0 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_98.vcd");
  if(my_type==0 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_99.vcd");
  if(my_type==0 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_100.vcd");
  if(my_type==0 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_101.vcd");
  if(my_type==0 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_102.vcd");
  if(my_type==0 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_103.vcd");
  if(my_type==0 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_104.vcd");
  if(my_type==0 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_105.vcd");
  if(my_type==0 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_106.vcd");
  if(my_type==0 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_107.vcd");
  if(my_type==0 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_108.vcd");
  if(my_type==0 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_109.vcd");
  if(my_type==0 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_110.vcd");
  if(my_type==0 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_111.vcd");
  if(my_type==0 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_112.vcd");
  if(my_type==0 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_113.vcd");
  if(my_type==0 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_114.vcd");
  if(my_type==0 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_115.vcd");
  if(my_type==0 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_116.vcd");
  if(my_type==0 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_117.vcd");
  if(my_type==0 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_118.vcd");
  if(my_type==0 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_119.vcd");
  if(my_type==0 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_120.vcd");
  if(my_type==0 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_121.vcd");
  if(my_type==0 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_122.vcd");
  if(my_type==0 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_123.vcd");
  if(my_type==0 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_124.vcd");
  if(my_type==0 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_125.vcd");
  if(my_type==0 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_126.vcd");
  if(my_type==0 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_127.vcd");
  if(my_type==0 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_128.vcd");
  if(my_type==0 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_129.vcd");
  if(my_type==0 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_130.vcd");
  if(my_type==0 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_131.vcd");
  if(my_type==0 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_132.vcd");
  if(my_type==0 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_133.vcd");
  if(my_type==0 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_134.vcd");
  if(my_type==0 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_135.vcd");
  if(my_type==0 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_136.vcd");
  if(my_type==0 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_137.vcd");
  if(my_type==0 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_138.vcd");
  if(my_type==0 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_139.vcd");
  if(my_type==0 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_140.vcd");
  if(my_type==0 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_141.vcd");
  if(my_type==0 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_142.vcd");
  if(my_type==0 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_143.vcd");
  if(my_type==0 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_144.vcd");
  if(my_type==0 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_145.vcd");
  if(my_type==0 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_146.vcd");
  if(my_type==0 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_147.vcd");
  if(my_type==0 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_148.vcd");
  if(my_type==0 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_149.vcd");
  if(my_type==0 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_150.vcd");
  if(my_type==0 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_151.vcd");
  if(my_type==0 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_152.vcd");
  if(my_type==0 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_153.vcd");
  if(my_type==0 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_154.vcd");
  if(my_type==0 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_155.vcd");
  if(my_type==0 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_156.vcd");
  if(my_type==0 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_157.vcd");
  if(my_type==0 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_158.vcd");
  if(my_type==0 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_159.vcd");
  if(my_type==0 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_160.vcd");
  if(my_type==0 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_161.vcd");
  if(my_type==0 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_162.vcd");
  if(my_type==0 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_163.vcd");
  if(my_type==0 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_164.vcd");
  if(my_type==0 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_165.vcd");
  if(my_type==0 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_166.vcd");
  if(my_type==0 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_167.vcd");
  if(my_type==0 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_168.vcd");
  if(my_type==0 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_169.vcd");
  if(my_type==0 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_170.vcd");
  if(my_type==0 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_171.vcd");
  if(my_type==0 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_172.vcd");
  if(my_type==0 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_173.vcd");
  if(my_type==0 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_174.vcd");
  if(my_type==0 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_175.vcd");
  if(my_type==0 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_176.vcd");
  if(my_type==0 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_177.vcd");
  if(my_type==0 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_178.vcd");
  if(my_type==0 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_179.vcd");
  if(my_type==0 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_180.vcd");
  if(my_type==0 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_181.vcd");
  if(my_type==0 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_182.vcd");
  if(my_type==0 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_183.vcd");
  if(my_type==0 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_184.vcd");
  if(my_type==0 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_185.vcd");
  if(my_type==0 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_186.vcd");
  if(my_type==0 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_187.vcd");
  if(my_type==0 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_188.vcd");
  if(my_type==0 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_189.vcd");
  if(my_type==0 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_190.vcd");
  if(my_type==0 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_191.vcd");
  if(my_type==0 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_192.vcd");
  if(my_type==0 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_193.vcd");
  if(my_type==0 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_194.vcd");
  if(my_type==0 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_195.vcd");
  if(my_type==0 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_196.vcd");
  if(my_type==0 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_197.vcd");
  if(my_type==0 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_198.vcd");
  if(my_type==0 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_199.vcd");
  if(my_type==0 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_200.vcd");
  if(my_type==0 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_201.vcd");
  if(my_type==0 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_202.vcd");
  if(my_type==0 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_203.vcd");
  if(my_type==0 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_204.vcd");
  if(my_type==0 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_205.vcd");
  if(my_type==0 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_206.vcd");
  if(my_type==0 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_207.vcd");
  if(my_type==0 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_208.vcd");
  if(my_type==0 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_209.vcd");
  if(my_type==0 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_210.vcd");
  if(my_type==0 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_211.vcd");
  if(my_type==0 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_212.vcd");
  if(my_type==0 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_213.vcd");
  if(my_type==0 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_214.vcd");
  if(my_type==0 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_215.vcd");
  if(my_type==0 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_216.vcd");
  if(my_type==0 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_217.vcd");
  if(my_type==0 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_218.vcd");
  if(my_type==0 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_219.vcd");
  if(my_type==0 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_220.vcd");
  if(my_type==0 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_221.vcd");
  if(my_type==0 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_222.vcd");
  if(my_type==0 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_223.vcd");
  if(my_type==0 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_224.vcd");
  if(my_type==0 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_225.vcd");
  if(my_type==0 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_226.vcd");
  if(my_type==0 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_227.vcd");
  if(my_type==0 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_228.vcd");
  if(my_type==0 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_229.vcd");
  if(my_type==0 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_230.vcd");
  if(my_type==0 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_231.vcd");
  if(my_type==0 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_232.vcd");
  if(my_type==0 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_233.vcd");
  if(my_type==0 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_234.vcd");
  if(my_type==0 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_235.vcd");
  if(my_type==0 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_236.vcd");
  if(my_type==0 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_237.vcd");
  if(my_type==0 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_238.vcd");
  if(my_type==0 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_239.vcd");
  if(my_type==0 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_240.vcd");
  if(my_type==0 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_241.vcd");
  if(my_type==0 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_242.vcd");
  if(my_type==0 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_243.vcd");
  if(my_type==0 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_244.vcd");
  if(my_type==0 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_245.vcd");
  if(my_type==0 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_246.vcd");
  if(my_type==0 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_247.vcd");
  if(my_type==0 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_248.vcd");
  if(my_type==0 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_249.vcd");
  if(my_type==0 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_250.vcd");
  if(my_type==0 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_251.vcd");
  if(my_type==0 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_252.vcd");
  if(my_type==0 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_253.vcd");
  if(my_type==0 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_254.vcd");
  if(my_type==0 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_255.vcd");
  if(my_type==0 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_256.vcd");
  if(my_type==0 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_257.vcd");
  if(my_type==0 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_258.vcd");
  if(my_type==0 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_259.vcd");
  if(my_type==0 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_260.vcd");
  if(my_type==0 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_261.vcd");
  if(my_type==0 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_262.vcd");
  if(my_type==0 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_263.vcd");
  if(my_type==0 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_264.vcd");
  if(my_type==0 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_265.vcd");
  if(my_type==0 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_266.vcd");
  if(my_type==0 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_267.vcd");
  if(my_type==0 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_268.vcd");
  if(my_type==0 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_269.vcd");
  if(my_type==0 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_270.vcd");
  if(my_type==0 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_271.vcd");
  if(my_type==0 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_272.vcd");
  if(my_type==0 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_273.vcd");
  if(my_type==0 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_274.vcd");
  if(my_type==0 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_275.vcd");
  if(my_type==0 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_276.vcd");
  if(my_type==0 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_277.vcd");
  if(my_type==0 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_278.vcd");
  if(my_type==0 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_279.vcd");
  if(my_type==0 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_280.vcd");
  if(my_type==0 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_281.vcd");
  if(my_type==0 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_282.vcd");
  if(my_type==0 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_283.vcd");
  if(my_type==0 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_284.vcd");
  if(my_type==0 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_285.vcd");
  if(my_type==0 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_286.vcd");
  if(my_type==0 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_287.vcd");
  if(my_type==0 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_288.vcd");
  if(my_type==0 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_289.vcd");
  if(my_type==0 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_290.vcd");
  if(my_type==0 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_291.vcd");
  if(my_type==0 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_292.vcd");
  if(my_type==0 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_293.vcd");
  if(my_type==0 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_294.vcd");
  if(my_type==0 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_295.vcd");
  if(my_type==0 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_296.vcd");
  if(my_type==0 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_297.vcd");
  if(my_type==0 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_298.vcd");
  if(my_type==0 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_299.vcd");
  if(my_type==0 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_300.vcd");
  if(my_type==0 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_301.vcd");
  if(my_type==0 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_302.vcd");
  if(my_type==0 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_303.vcd");
  if(my_type==0 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_304.vcd");
  if(my_type==0 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_305.vcd");
  if(my_type==0 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_306.vcd");
  if(my_type==0 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_307.vcd");
  if(my_type==0 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_308.vcd");
  if(my_type==0 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_309.vcd");
  if(my_type==0 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_310.vcd");
  if(my_type==0 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_311.vcd");
  if(my_type==0 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_312.vcd");
  if(my_type==0 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_313.vcd");
  if(my_type==0 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_314.vcd");
  if(my_type==0 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_315.vcd");
  if(my_type==0 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_316.vcd");
  if(my_type==0 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_317.vcd");
  if(my_type==0 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_318.vcd");
  if(my_type==0 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_319.vcd");
  if(my_type==0 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_320.vcd");
  if(my_type==0 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_321.vcd");
  if(my_type==0 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_322.vcd");
  if(my_type==0 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_323.vcd");
  if(my_type==0 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_324.vcd");
  if(my_type==0 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_325.vcd");
  if(my_type==0 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_326.vcd");
  if(my_type==0 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_327.vcd");
  if(my_type==0 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_328.vcd");
  if(my_type==0 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_329.vcd");
  if(my_type==0 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_330.vcd");
  if(my_type==0 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_331.vcd");
  if(my_type==0 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_332.vcd");
  if(my_type==0 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_333.vcd");
  if(my_type==0 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_334.vcd");
  if(my_type==0 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_335.vcd");
  if(my_type==0 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_336.vcd");
  if(my_type==0 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_337.vcd");
  if(my_type==0 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_338.vcd");
  if(my_type==0 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_339.vcd");
  if(my_type==0 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_340.vcd");
  if(my_type==0 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_341.vcd");
  if(my_type==0 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_342.vcd");
  if(my_type==0 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_343.vcd");
  if(my_type==0 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_344.vcd");
  if(my_type==0 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_345.vcd");
  if(my_type==0 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_346.vcd");
  if(my_type==0 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_347.vcd");
  if(my_type==0 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_348.vcd");
  if(my_type==0 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_349.vcd");
  if(my_type==0 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_350.vcd");
  if(my_type==0 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_351.vcd");
  if(my_type==0 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_352.vcd");
  if(my_type==0 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_353.vcd");
  if(my_type==0 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_354.vcd");
  if(my_type==0 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_355.vcd");
  if(my_type==0 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_356.vcd");
  if(my_type==0 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_357.vcd");
  if(my_type==0 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_358.vcd");
  if(my_type==0 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_359.vcd");
  if(my_type==0 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_360.vcd");
  if(my_type==0 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_361.vcd");
  if(my_type==0 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_362.vcd");
  if(my_type==0 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_363.vcd");
  if(my_type==0 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_364.vcd");
  if(my_type==0 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_365.vcd");
  if(my_type==0 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_366.vcd");
  if(my_type==0 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_367.vcd");
  if(my_type==0 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_368.vcd");
  if(my_type==0 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_369.vcd");
  if(my_type==0 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_370.vcd");
  if(my_type==0 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_371.vcd");
  if(my_type==0 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_372.vcd");
  if(my_type==0 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_373.vcd");
  if(my_type==0 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_374.vcd");
  if(my_type==0 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_375.vcd");
  if(my_type==0 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_376.vcd");
  if(my_type==0 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_377.vcd");
  if(my_type==0 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_378.vcd");
  if(my_type==0 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_379.vcd");
  if(my_type==0 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_380.vcd");
  if(my_type==0 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_381.vcd");
  if(my_type==0 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_382.vcd");
  if(my_type==0 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_383.vcd");
  if(my_type==0 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_384.vcd");
  if(my_type==0 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_385.vcd");
  if(my_type==0 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_386.vcd");
  if(my_type==0 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_387.vcd");
  if(my_type==0 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_388.vcd");
  if(my_type==0 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_389.vcd");
  if(my_type==0 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_390.vcd");
  if(my_type==0 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_391.vcd");
  if(my_type==0 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_392.vcd");
  if(my_type==0 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_393.vcd");
  if(my_type==0 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_394.vcd");
  if(my_type==0 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_395.vcd");
  if(my_type==0 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_396.vcd");
  if(my_type==0 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_397.vcd");
  if(my_type==0 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_398.vcd");
  if(my_type==0 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_399.vcd");
  if(my_type==0 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_400.vcd");
  if(my_type==0 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_401.vcd");
  if(my_type==0 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_402.vcd");
  if(my_type==0 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_403.vcd");
  if(my_type==0 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_404.vcd");
  if(my_type==0 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_405.vcd");
  if(my_type==0 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_406.vcd");
  if(my_type==0 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_407.vcd");
  if(my_type==0 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_408.vcd");
  if(my_type==0 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_409.vcd");
  if(my_type==0 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_410.vcd");
  if(my_type==0 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_411.vcd");
  if(my_type==0 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_412.vcd");
  if(my_type==0 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_413.vcd");
  if(my_type==0 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_414.vcd");
  if(my_type==0 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_415.vcd");
  if(my_type==0 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_416.vcd");
  if(my_type==0 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_417.vcd");
  if(my_type==0 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_418.vcd");
  if(my_type==0 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_419.vcd");
  if(my_type==0 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_420.vcd");
  if(my_type==0 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_421.vcd");
  if(my_type==0 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_422.vcd");
  if(my_type==0 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_423.vcd");
  if(my_type==0 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_424.vcd");
  if(my_type==0 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_425.vcd");
  if(my_type==0 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_426.vcd");
  if(my_type==0 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_427.vcd");
  if(my_type==0 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_428.vcd");
  if(my_type==0 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_429.vcd");
  if(my_type==0 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_430.vcd");
  if(my_type==0 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_431.vcd");
  if(my_type==0 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_432.vcd");
  if(my_type==0 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_433.vcd");
  if(my_type==0 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_434.vcd");
  if(my_type==0 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_435.vcd");
  if(my_type==0 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_436.vcd");
  if(my_type==0 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_437.vcd");
  if(my_type==0 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_438.vcd");
  if(my_type==0 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_439.vcd");
  if(my_type==0 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_440.vcd");
  if(my_type==0 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_441.vcd");
  if(my_type==0 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_442.vcd");
  if(my_type==0 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_443.vcd");
  if(my_type==0 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_444.vcd");
  if(my_type==0 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_445.vcd");
  if(my_type==0 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_446.vcd");
  if(my_type==0 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_447.vcd");
  if(my_type==0 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_448.vcd");
  if(my_type==0 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_449.vcd");
  if(my_type==0 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_450.vcd");
  if(my_type==0 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_451.vcd");
  if(my_type==0 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_452.vcd");
  if(my_type==0 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_453.vcd");
  if(my_type==0 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_454.vcd");
  if(my_type==0 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_455.vcd");
  if(my_type==0 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_456.vcd");
  if(my_type==0 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_457.vcd");
  if(my_type==0 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_458.vcd");
  if(my_type==0 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_459.vcd");
  if(my_type==0 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_460.vcd");
  if(my_type==0 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_461.vcd");
  if(my_type==0 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_462.vcd");
  if(my_type==0 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_463.vcd");
  if(my_type==0 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_464.vcd");
  if(my_type==0 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_465.vcd");
  if(my_type==0 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_466.vcd");
  if(my_type==0 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_467.vcd");
  if(my_type==0 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_468.vcd");
  if(my_type==0 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_469.vcd");
  if(my_type==0 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_470.vcd");
  if(my_type==0 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_471.vcd");
  if(my_type==0 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_472.vcd");
  if(my_type==0 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_473.vcd");
  if(my_type==0 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_474.vcd");
  if(my_type==0 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_475.vcd");
  if(my_type==0 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_476.vcd");
  if(my_type==0 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_477.vcd");
  if(my_type==0 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_478.vcd");
  if(my_type==0 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_479.vcd");
  if(my_type==0 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_480.vcd");
  if(my_type==0 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_481.vcd");
  if(my_type==0 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_482.vcd");
  if(my_type==0 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_483.vcd");
  if(my_type==0 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_484.vcd");
  if(my_type==0 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_485.vcd");
  if(my_type==0 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_486.vcd");
  if(my_type==0 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_487.vcd");
  if(my_type==0 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_488.vcd");
  if(my_type==0 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_489.vcd");
  if(my_type==0 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_490.vcd");
  if(my_type==0 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_491.vcd");
  if(my_type==0 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_492.vcd");
  if(my_type==0 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_493.vcd");
  if(my_type==0 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_494.vcd");
  if(my_type==0 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_495.vcd");
  if(my_type==0 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_496.vcd");
  if(my_type==0 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_497.vcd");
  if(my_type==0 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_498.vcd");
  if(my_type==0 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_499.vcd");
  if(my_type==0 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_500.vcd");
  if(my_type==0 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_501.vcd");
  if(my_type==0 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_502.vcd");
  if(my_type==0 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_503.vcd");
  if(my_type==0 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_504.vcd");
  if(my_type==0 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_505.vcd");
  if(my_type==0 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_506.vcd");
  if(my_type==0 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_507.vcd");
  if(my_type==0 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_508.vcd");
  if(my_type==0 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_509.vcd");
  if(my_type==0 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_510.vcd");
  if(my_type==0 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_511.vcd");
  if(my_type==0 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_512.vcd");
  if(my_type==0 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_513.vcd");
  if(my_type==0 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_514.vcd");
  if(my_type==0 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_515.vcd");
  if(my_type==0 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_516.vcd");
  if(my_type==0 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_517.vcd");
  if(my_type==0 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_518.vcd");
  if(my_type==0 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_519.vcd");
  if(my_type==0 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_520.vcd");
  if(my_type==0 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_521.vcd");
  if(my_type==0 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_522.vcd");
  if(my_type==0 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_523.vcd");
  if(my_type==0 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_524.vcd");
  if(my_type==0 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_525.vcd");
  if(my_type==0 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_526.vcd");
  if(my_type==0 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_527.vcd");
  if(my_type==0 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_528.vcd");
  if(my_type==0 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_529.vcd");
  if(my_type==0 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_530.vcd");
  if(my_type==0 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_531.vcd");
  if(my_type==0 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_532.vcd");
  if(my_type==0 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_533.vcd");
  if(my_type==0 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_534.vcd");
  if(my_type==0 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_535.vcd");
  if(my_type==0 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_536.vcd");
  if(my_type==0 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_537.vcd");
  if(my_type==0 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_538.vcd");
  if(my_type==0 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_539.vcd");
  if(my_type==0 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_540.vcd");
  if(my_type==0 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_541.vcd");
  if(my_type==0 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_542.vcd");
  if(my_type==0 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_543.vcd");
  if(my_type==0 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_544.vcd");
  if(my_type==0 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_545.vcd");
  if(my_type==0 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_546.vcd");
  if(my_type==0 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_547.vcd");
  if(my_type==0 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_548.vcd");
  if(my_type==0 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_549.vcd");
  if(my_type==0 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_550.vcd");
  if(my_type==0 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_551.vcd");
  if(my_type==0 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_552.vcd");
  if(my_type==0 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_553.vcd");
  if(my_type==0 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_554.vcd");
  if(my_type==0 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_555.vcd");
  if(my_type==0 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_556.vcd");
  if(my_type==0 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_557.vcd");
  if(my_type==0 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_558.vcd");
  if(my_type==0 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_559.vcd");
  if(my_type==0 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_560.vcd");
  if(my_type==0 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_561.vcd");
  if(my_type==0 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_562.vcd");
  if(my_type==0 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_563.vcd");
  if(my_type==0 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_564.vcd");
  if(my_type==0 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_565.vcd");
  if(my_type==0 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_566.vcd");
  if(my_type==0 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_567.vcd");
  if(my_type==0 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_568.vcd");
  if(my_type==0 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_569.vcd");
  if(my_type==0 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_570.vcd");
  if(my_type==0 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_571.vcd");
  if(my_type==0 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_572.vcd");
  if(my_type==0 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_573.vcd");
  if(my_type==0 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_574.vcd");
  if(my_type==0 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_575.vcd");
  if(my_type==0 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_576.vcd");
  if(my_type==0 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_577.vcd");
  if(my_type==0 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_578.vcd");
  if(my_type==0 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_579.vcd");
  if(my_type==0 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_580.vcd");
  if(my_type==0 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_581.vcd");
  if(my_type==0 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_582.vcd");
  if(my_type==0 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_583.vcd");
  if(my_type==0 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_584.vcd");
  if(my_type==0 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_585.vcd");
  if(my_type==0 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_586.vcd");
  if(my_type==0 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_587.vcd");
  if(my_type==0 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_588.vcd");
  if(my_type==0 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_589.vcd");
  if(my_type==0 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_590.vcd");
  if(my_type==0 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_591.vcd");
  if(my_type==0 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_592.vcd");
  if(my_type==0 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_593.vcd");
  if(my_type==0 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_594.vcd");
  if(my_type==0 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_595.vcd");
  if(my_type==0 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_596.vcd");
  if(my_type==0 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_597.vcd");
  if(my_type==0 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_598.vcd");
  if(my_type==0 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_599.vcd");
  if(my_type==0 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_600.vcd");
  if(my_type==0 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_601.vcd");
  if(my_type==0 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_602.vcd");
  if(my_type==0 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_603.vcd");
  if(my_type==0 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_604.vcd");
  if(my_type==0 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_605.vcd");
  if(my_type==0 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_606.vcd");
  if(my_type==0 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_607.vcd");
  if(my_type==0 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_608.vcd");
  if(my_type==0 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_609.vcd");
  if(my_type==0 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_610.vcd");
  if(my_type==0 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_611.vcd");
  if(my_type==0 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_612.vcd");
  if(my_type==0 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_613.vcd");
  if(my_type==0 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_614.vcd");
  if(my_type==0 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_615.vcd");
  if(my_type==0 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_616.vcd");
  if(my_type==0 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_617.vcd");
  if(my_type==0 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_618.vcd");
  if(my_type==0 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_619.vcd");
  if(my_type==0 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_620.vcd");
  if(my_type==0 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_621.vcd");
  if(my_type==0 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_622.vcd");
  if(my_type==0 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_623.vcd");
  if(my_type==0 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_624.vcd");
  if(my_type==0 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_625.vcd");
  if(my_type==0 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_626.vcd");
  if(my_type==0 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_627.vcd");
  if(my_type==0 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_628.vcd");
  if(my_type==0 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_629.vcd");
  if(my_type==0 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_630.vcd");
  if(my_type==0 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_631.vcd");
  if(my_type==0 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_632.vcd");
  if(my_type==0 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_633.vcd");
  if(my_type==0 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_634.vcd");
  if(my_type==0 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_635.vcd");
  if(my_type==0 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_636.vcd");
  if(my_type==0 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_637.vcd");
  if(my_type==0 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_638.vcd");
  if(my_type==0 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_639.vcd");
  if(my_type==0 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_640.vcd");
  if(my_type==0 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_641.vcd");
  if(my_type==0 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_642.vcd");
  if(my_type==0 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_643.vcd");
  if(my_type==0 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_644.vcd");
  if(my_type==0 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_645.vcd");
  if(my_type==0 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_646.vcd");
  if(my_type==0 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_647.vcd");
  if(my_type==0 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_648.vcd");
  if(my_type==0 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_649.vcd");
  if(my_type==0 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_650.vcd");
  if(my_type==0 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_651.vcd");
  if(my_type==0 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_652.vcd");
  if(my_type==0 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_653.vcd");
  if(my_type==0 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_654.vcd");
  if(my_type==0 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_655.vcd");
  if(my_type==0 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_656.vcd");
  if(my_type==0 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_657.vcd");
  if(my_type==0 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_658.vcd");
  if(my_type==0 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_659.vcd");
  if(my_type==0 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_660.vcd");
  if(my_type==0 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_661.vcd");
  if(my_type==0 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_662.vcd");
  if(my_type==0 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_663.vcd");
  if(my_type==0 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_664.vcd");
  if(my_type==0 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_665.vcd");
  if(my_type==0 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_666.vcd");
  if(my_type==0 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_667.vcd");
  if(my_type==0 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_668.vcd");
  if(my_type==0 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_669.vcd");
  if(my_type==0 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_670.vcd");
  if(my_type==0 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_671.vcd");
  if(my_type==0 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_672.vcd");
  if(my_type==0 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_673.vcd");
  if(my_type==0 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_674.vcd");
  if(my_type==0 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_675.vcd");
  if(my_type==0 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_676.vcd");
  if(my_type==0 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_677.vcd");
  if(my_type==0 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_678.vcd");
  if(my_type==0 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_679.vcd");
  if(my_type==0 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_680.vcd");
  if(my_type==0 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_681.vcd");
  if(my_type==0 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_682.vcd");
  if(my_type==0 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_683.vcd");
  if(my_type==0 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_684.vcd");
  if(my_type==0 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_685.vcd");
  if(my_type==0 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_686.vcd");
  if(my_type==0 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_687.vcd");
  if(my_type==0 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_688.vcd");
  if(my_type==0 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_689.vcd");
  if(my_type==0 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_690.vcd");
  if(my_type==0 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_691.vcd");
  if(my_type==0 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_692.vcd");
  if(my_type==0 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_693.vcd");
  if(my_type==0 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_694.vcd");
  if(my_type==0 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_695.vcd");
  if(my_type==0 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_696.vcd");
  if(my_type==0 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_697.vcd");
  if(my_type==0 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_698.vcd");
  if(my_type==0 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_699.vcd");
  if(my_type==0 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_700.vcd");
  if(my_type==0 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_701.vcd");
  if(my_type==0 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_702.vcd");
  if(my_type==0 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_703.vcd");
  if(my_type==0 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_704.vcd");
  if(my_type==0 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_705.vcd");
  if(my_type==0 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_706.vcd");
  if(my_type==0 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_707.vcd");
  if(my_type==0 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_708.vcd");
  if(my_type==0 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_709.vcd");
  if(my_type==0 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_710.vcd");
  if(my_type==0 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_711.vcd");
  if(my_type==0 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_712.vcd");
  if(my_type==0 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_713.vcd");
  if(my_type==0 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_714.vcd");
  if(my_type==0 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_715.vcd");
  if(my_type==0 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_716.vcd");
  if(my_type==0 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_717.vcd");
  if(my_type==0 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_718.vcd");
  if(my_type==0 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_719.vcd");
  if(my_type==0 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_720.vcd");
  if(my_type==0 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_721.vcd");
  if(my_type==0 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_722.vcd");
  if(my_type==0 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_723.vcd");
  if(my_type==0 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_724.vcd");
  if(my_type==0 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_725.vcd");
  if(my_type==0 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_726.vcd");
  if(my_type==0 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_727.vcd");
  if(my_type==0 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_728.vcd");
  if(my_type==0 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_729.vcd");
  if(my_type==0 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_730.vcd");
  if(my_type==0 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_731.vcd");
  if(my_type==0 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_732.vcd");
  if(my_type==0 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_733.vcd");
  if(my_type==0 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_734.vcd");
  if(my_type==0 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_735.vcd");
  if(my_type==0 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_736.vcd");
  if(my_type==0 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_737.vcd");
  if(my_type==0 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_738.vcd");
  if(my_type==0 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_739.vcd");
  if(my_type==0 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_740.vcd");
  if(my_type==0 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_741.vcd");
  if(my_type==0 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_742.vcd");
  if(my_type==0 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_743.vcd");
  if(my_type==0 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_744.vcd");
  if(my_type==0 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_745.vcd");
  if(my_type==0 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_746.vcd");
  if(my_type==0 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_747.vcd");
  if(my_type==0 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_748.vcd");
  if(my_type==0 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_749.vcd");
  if(my_type==0 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_750.vcd");
  if(my_type==0 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_751.vcd");
  if(my_type==0 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_752.vcd");
  if(my_type==0 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_753.vcd");
  if(my_type==0 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_754.vcd");
  if(my_type==0 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_755.vcd");
  if(my_type==0 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_756.vcd");
  if(my_type==0 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_757.vcd");
  if(my_type==0 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_758.vcd");
  if(my_type==0 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_759.vcd");
  if(my_type==0 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_760.vcd");
  if(my_type==0 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_761.vcd");
  if(my_type==0 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_762.vcd");
  if(my_type==0 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_763.vcd");
  if(my_type==0 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_764.vcd");
  if(my_type==0 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_765.vcd");
  if(my_type==0 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_766.vcd");
  if(my_type==0 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_767.vcd");
  if(my_type==0 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_768.vcd");
  if(my_type==0 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_769.vcd");
  if(my_type==0 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_770.vcd");
  if(my_type==0 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_771.vcd");
  if(my_type==0 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_772.vcd");
  if(my_type==0 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_773.vcd");
  if(my_type==0 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_774.vcd");
  if(my_type==0 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_775.vcd");
  if(my_type==0 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_776.vcd");
  if(my_type==0 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_777.vcd");
  if(my_type==0 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_778.vcd");
  if(my_type==0 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_779.vcd");
  if(my_type==0 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_780.vcd");
  if(my_type==0 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_781.vcd");
  if(my_type==0 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_782.vcd");
  if(my_type==0 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_783.vcd");
  if(my_type==0 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_784.vcd");
  if(my_type==0 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_785.vcd");
  if(my_type==0 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_786.vcd");
  if(my_type==0 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_787.vcd");
  if(my_type==0 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_788.vcd");
  if(my_type==0 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_789.vcd");
  if(my_type==0 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_790.vcd");
  if(my_type==0 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_791.vcd");
  if(my_type==0 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_792.vcd");
  if(my_type==0 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_793.vcd");
  if(my_type==0 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_794.vcd");
  if(my_type==0 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_795.vcd");
  if(my_type==0 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_796.vcd");
  if(my_type==0 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_797.vcd");
  if(my_type==0 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_798.vcd");
  if(my_type==0 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_799.vcd");
  if(my_type==0 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_800.vcd");
  if(my_type==0 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_801.vcd");
  if(my_type==0 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_802.vcd");
  if(my_type==0 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_803.vcd");
  if(my_type==0 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_804.vcd");
  if(my_type==0 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_805.vcd");
  if(my_type==0 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_806.vcd");
  if(my_type==0 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_807.vcd");
  if(my_type==0 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_808.vcd");
  if(my_type==0 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_809.vcd");
  if(my_type==0 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_810.vcd");
  if(my_type==0 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_811.vcd");
  if(my_type==0 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_812.vcd");
  if(my_type==0 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_813.vcd");
  if(my_type==0 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_814.vcd");
  if(my_type==0 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_815.vcd");
  if(my_type==0 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_816.vcd");
  if(my_type==0 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_817.vcd");
  if(my_type==0 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_818.vcd");
  if(my_type==0 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_819.vcd");
  if(my_type==0 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_820.vcd");
  if(my_type==0 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_821.vcd");
  if(my_type==0 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_822.vcd");
  if(my_type==0 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_823.vcd");
  if(my_type==0 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_824.vcd");
  if(my_type==0 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_825.vcd");
  if(my_type==0 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_826.vcd");
  if(my_type==0 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_827.vcd");
  if(my_type==0 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_828.vcd");
  if(my_type==0 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_829.vcd");
  if(my_type==0 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_830.vcd");
  if(my_type==0 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_831.vcd");
  if(my_type==0 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_832.vcd");
  if(my_type==0 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_833.vcd");
  if(my_type==0 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_834.vcd");
  if(my_type==0 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_835.vcd");
  if(my_type==0 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_836.vcd");
  if(my_type==0 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_837.vcd");
  if(my_type==0 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_838.vcd");
  if(my_type==0 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_839.vcd");
  if(my_type==0 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_840.vcd");
  if(my_type==0 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_841.vcd");
  if(my_type==0 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_842.vcd");
  if(my_type==0 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_843.vcd");
  if(my_type==0 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_844.vcd");
  if(my_type==0 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_845.vcd");
  if(my_type==0 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_846.vcd");
  if(my_type==0 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_847.vcd");
  if(my_type==0 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_848.vcd");
  if(my_type==0 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_849.vcd");
  if(my_type==0 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_850.vcd");
  if(my_type==0 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_851.vcd");
  if(my_type==0 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_852.vcd");
  if(my_type==0 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_853.vcd");
  if(my_type==0 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_854.vcd");
  if(my_type==0 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_855.vcd");
  if(my_type==0 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_856.vcd");
  if(my_type==0 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_857.vcd");
  if(my_type==0 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_858.vcd");
  if(my_type==0 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_859.vcd");
  if(my_type==0 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_860.vcd");
  if(my_type==0 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_861.vcd");
  if(my_type==0 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_862.vcd");
  if(my_type==0 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_863.vcd");
  if(my_type==0 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_864.vcd");
  if(my_type==0 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_865.vcd");
  if(my_type==0 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_866.vcd");
  if(my_type==0 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_867.vcd");
  if(my_type==0 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_868.vcd");
  if(my_type==0 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_869.vcd");
  if(my_type==0 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_870.vcd");
  if(my_type==0 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_871.vcd");
  if(my_type==0 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_872.vcd");
  if(my_type==0 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_873.vcd");
  if(my_type==0 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_874.vcd");
  if(my_type==0 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_875.vcd");
  if(my_type==0 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_876.vcd");
  if(my_type==0 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_877.vcd");
  if(my_type==0 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_878.vcd");
  if(my_type==0 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_879.vcd");
  if(my_type==0 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_880.vcd");
  if(my_type==0 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_881.vcd");
  if(my_type==0 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_882.vcd");
  if(my_type==0 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_883.vcd");
  if(my_type==0 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_884.vcd");
  if(my_type==0 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_885.vcd");
  if(my_type==0 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_886.vcd");
  if(my_type==0 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_887.vcd");
  if(my_type==0 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_888.vcd");
  if(my_type==0 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_889.vcd");
  if(my_type==0 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_890.vcd");
  if(my_type==0 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_891.vcd");
  if(my_type==0 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_892.vcd");
  if(my_type==0 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_893.vcd");
  if(my_type==0 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_894.vcd");
  if(my_type==0 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_895.vcd");
  if(my_type==0 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_896.vcd");
  if(my_type==0 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_897.vcd");
  if(my_type==0 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_898.vcd");
  if(my_type==0 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_899.vcd");
  if(my_type==0 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_900.vcd");
  if(my_type==0 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_901.vcd");
  if(my_type==0 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_902.vcd");
  if(my_type==0 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_903.vcd");
  if(my_type==0 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_904.vcd");
  if(my_type==0 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_905.vcd");
  if(my_type==0 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_906.vcd");
  if(my_type==0 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_907.vcd");
  if(my_type==0 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_908.vcd");
  if(my_type==0 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_909.vcd");
  if(my_type==0 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_910.vcd");
  if(my_type==0 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_911.vcd");
  if(my_type==0 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_912.vcd");
  if(my_type==0 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_913.vcd");
  if(my_type==0 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_914.vcd");
  if(my_type==0 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_915.vcd");
  if(my_type==0 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_916.vcd");
  if(my_type==0 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_917.vcd");
  if(my_type==0 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_918.vcd");
  if(my_type==0 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_919.vcd");
  if(my_type==0 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_920.vcd");
  if(my_type==0 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_921.vcd");
  if(my_type==0 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_922.vcd");
  if(my_type==0 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_923.vcd");
  if(my_type==0 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_924.vcd");
  if(my_type==0 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_925.vcd");
  if(my_type==0 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_926.vcd");
  if(my_type==0 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_927.vcd");
  if(my_type==0 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_928.vcd");
  if(my_type==0 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_929.vcd");
  if(my_type==0 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_930.vcd");
  if(my_type==0 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_931.vcd");
  if(my_type==0 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_932.vcd");
  if(my_type==0 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_933.vcd");
  if(my_type==0 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_934.vcd");
  if(my_type==0 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_935.vcd");
  if(my_type==0 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_936.vcd");
  if(my_type==0 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_937.vcd");
  if(my_type==0 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_938.vcd");
  if(my_type==0 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_939.vcd");
  if(my_type==0 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_940.vcd");
  if(my_type==0 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_941.vcd");
  if(my_type==0 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_942.vcd");
  if(my_type==0 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_943.vcd");
  if(my_type==0 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_944.vcd");
  if(my_type==0 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_945.vcd");
  if(my_type==0 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_946.vcd");
  if(my_type==0 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_947.vcd");
  if(my_type==0 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_948.vcd");
  if(my_type==0 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_949.vcd");
  if(my_type==0 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_950.vcd");
  if(my_type==0 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_951.vcd");
  if(my_type==0 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_952.vcd");
  if(my_type==0 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_953.vcd");
  if(my_type==0 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_954.vcd");
  if(my_type==0 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_955.vcd");
  if(my_type==0 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_956.vcd");
  if(my_type==0 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_957.vcd");
  if(my_type==0 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_958.vcd");
  if(my_type==0 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_959.vcd");
  if(my_type==0 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_960.vcd");
  if(my_type==0 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_961.vcd");
  if(my_type==0 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_962.vcd");
  if(my_type==0 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_963.vcd");
  if(my_type==0 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_964.vcd");
  if(my_type==0 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_965.vcd");
  if(my_type==0 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_966.vcd");
  if(my_type==0 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_967.vcd");
  if(my_type==0 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_968.vcd");
  if(my_type==0 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_969.vcd");
  if(my_type==0 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_970.vcd");
  if(my_type==0 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_971.vcd");
  if(my_type==0 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_972.vcd");
  if(my_type==0 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_973.vcd");
  if(my_type==0 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_974.vcd");
  if(my_type==0 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_975.vcd");
  if(my_type==0 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_976.vcd");
  if(my_type==0 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_977.vcd");
  if(my_type==0 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_978.vcd");
  if(my_type==0 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_979.vcd");
  if(my_type==0 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_980.vcd");
  if(my_type==0 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_981.vcd");
  if(my_type==0 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_982.vcd");
  if(my_type==0 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_983.vcd");
  if(my_type==0 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_984.vcd");
  if(my_type==0 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_985.vcd");
  if(my_type==0 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_986.vcd");
  if(my_type==0 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_987.vcd");
  if(my_type==0 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_988.vcd");
  if(my_type==0 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_989.vcd");
  if(my_type==0 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_990.vcd");
  if(my_type==0 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_991.vcd");
  if(my_type==0 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_992.vcd");
  if(my_type==0 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_993.vcd");
  if(my_type==0 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_994.vcd");
  if(my_type==0 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_995.vcd");
  if(my_type==0 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_996.vcd");
  if(my_type==0 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_997.vcd");
  if(my_type==0 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_998.vcd");
  if(my_type==0 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_0_999.vcd");
  if(my_type==1 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_0.vcd");
  if(my_type==1 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_1.vcd");
  if(my_type==1 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_2.vcd");
  if(my_type==1 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_3.vcd");
  if(my_type==1 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_4.vcd");
  if(my_type==1 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_5.vcd");
  if(my_type==1 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_6.vcd");
  if(my_type==1 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_7.vcd");
  if(my_type==1 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_8.vcd");
  if(my_type==1 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_9.vcd");
  if(my_type==1 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_10.vcd");
  if(my_type==1 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_11.vcd");
  if(my_type==1 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_12.vcd");
  if(my_type==1 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_13.vcd");
  if(my_type==1 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_14.vcd");
  if(my_type==1 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_15.vcd");
  if(my_type==1 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_16.vcd");
  if(my_type==1 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_17.vcd");
  if(my_type==1 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_18.vcd");
  if(my_type==1 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_19.vcd");
  if(my_type==1 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_20.vcd");
  if(my_type==1 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_21.vcd");
  if(my_type==1 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_22.vcd");
  if(my_type==1 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_23.vcd");
  if(my_type==1 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_24.vcd");
  if(my_type==1 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_25.vcd");
  if(my_type==1 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_26.vcd");
  if(my_type==1 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_27.vcd");
  if(my_type==1 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_28.vcd");
  if(my_type==1 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_29.vcd");
  if(my_type==1 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_30.vcd");
  if(my_type==1 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_31.vcd");
  if(my_type==1 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_32.vcd");
  if(my_type==1 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_33.vcd");
  if(my_type==1 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_34.vcd");
  if(my_type==1 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_35.vcd");
  if(my_type==1 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_36.vcd");
  if(my_type==1 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_37.vcd");
  if(my_type==1 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_38.vcd");
  if(my_type==1 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_39.vcd");
  if(my_type==1 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_40.vcd");
  if(my_type==1 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_41.vcd");
  if(my_type==1 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_42.vcd");
  if(my_type==1 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_43.vcd");
  if(my_type==1 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_44.vcd");
  if(my_type==1 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_45.vcd");
  if(my_type==1 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_46.vcd");
  if(my_type==1 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_47.vcd");
  if(my_type==1 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_48.vcd");
  if(my_type==1 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_49.vcd");
  if(my_type==1 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_50.vcd");
  if(my_type==1 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_51.vcd");
  if(my_type==1 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_52.vcd");
  if(my_type==1 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_53.vcd");
  if(my_type==1 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_54.vcd");
  if(my_type==1 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_55.vcd");
  if(my_type==1 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_56.vcd");
  if(my_type==1 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_57.vcd");
  if(my_type==1 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_58.vcd");
  if(my_type==1 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_59.vcd");
  if(my_type==1 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_60.vcd");
  if(my_type==1 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_61.vcd");
  if(my_type==1 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_62.vcd");
  if(my_type==1 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_63.vcd");
  if(my_type==1 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_64.vcd");
  if(my_type==1 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_65.vcd");
  if(my_type==1 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_66.vcd");
  if(my_type==1 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_67.vcd");
  if(my_type==1 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_68.vcd");
  if(my_type==1 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_69.vcd");
  if(my_type==1 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_70.vcd");
  if(my_type==1 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_71.vcd");
  if(my_type==1 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_72.vcd");
  if(my_type==1 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_73.vcd");
  if(my_type==1 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_74.vcd");
  if(my_type==1 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_75.vcd");
  if(my_type==1 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_76.vcd");
  if(my_type==1 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_77.vcd");
  if(my_type==1 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_78.vcd");
  if(my_type==1 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_79.vcd");
  if(my_type==1 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_80.vcd");
  if(my_type==1 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_81.vcd");
  if(my_type==1 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_82.vcd");
  if(my_type==1 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_83.vcd");
  if(my_type==1 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_84.vcd");
  if(my_type==1 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_85.vcd");
  if(my_type==1 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_86.vcd");
  if(my_type==1 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_87.vcd");
  if(my_type==1 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_88.vcd");
  if(my_type==1 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_89.vcd");
  if(my_type==1 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_90.vcd");
  if(my_type==1 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_91.vcd");
  if(my_type==1 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_92.vcd");
  if(my_type==1 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_93.vcd");
  if(my_type==1 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_94.vcd");
  if(my_type==1 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_95.vcd");
  if(my_type==1 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_96.vcd");
  if(my_type==1 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_97.vcd");
  if(my_type==1 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_98.vcd");
  if(my_type==1 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_99.vcd");
  if(my_type==1 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_100.vcd");
  if(my_type==1 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_101.vcd");
  if(my_type==1 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_102.vcd");
  if(my_type==1 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_103.vcd");
  if(my_type==1 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_104.vcd");
  if(my_type==1 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_105.vcd");
  if(my_type==1 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_106.vcd");
  if(my_type==1 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_107.vcd");
  if(my_type==1 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_108.vcd");
  if(my_type==1 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_109.vcd");
  if(my_type==1 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_110.vcd");
  if(my_type==1 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_111.vcd");
  if(my_type==1 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_112.vcd");
  if(my_type==1 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_113.vcd");
  if(my_type==1 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_114.vcd");
  if(my_type==1 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_115.vcd");
  if(my_type==1 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_116.vcd");
  if(my_type==1 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_117.vcd");
  if(my_type==1 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_118.vcd");
  if(my_type==1 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_119.vcd");
  if(my_type==1 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_120.vcd");
  if(my_type==1 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_121.vcd");
  if(my_type==1 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_122.vcd");
  if(my_type==1 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_123.vcd");
  if(my_type==1 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_124.vcd");
  if(my_type==1 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_125.vcd");
  if(my_type==1 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_126.vcd");
  if(my_type==1 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_127.vcd");
  if(my_type==1 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_128.vcd");
  if(my_type==1 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_129.vcd");
  if(my_type==1 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_130.vcd");
  if(my_type==1 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_131.vcd");
  if(my_type==1 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_132.vcd");
  if(my_type==1 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_133.vcd");
  if(my_type==1 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_134.vcd");
  if(my_type==1 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_135.vcd");
  if(my_type==1 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_136.vcd");
  if(my_type==1 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_137.vcd");
  if(my_type==1 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_138.vcd");
  if(my_type==1 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_139.vcd");
  if(my_type==1 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_140.vcd");
  if(my_type==1 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_141.vcd");
  if(my_type==1 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_142.vcd");
  if(my_type==1 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_143.vcd");
  if(my_type==1 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_144.vcd");
  if(my_type==1 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_145.vcd");
  if(my_type==1 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_146.vcd");
  if(my_type==1 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_147.vcd");
  if(my_type==1 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_148.vcd");
  if(my_type==1 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_149.vcd");
  if(my_type==1 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_150.vcd");
  if(my_type==1 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_151.vcd");
  if(my_type==1 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_152.vcd");
  if(my_type==1 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_153.vcd");
  if(my_type==1 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_154.vcd");
  if(my_type==1 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_155.vcd");
  if(my_type==1 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_156.vcd");
  if(my_type==1 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_157.vcd");
  if(my_type==1 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_158.vcd");
  if(my_type==1 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_159.vcd");
  if(my_type==1 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_160.vcd");
  if(my_type==1 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_161.vcd");
  if(my_type==1 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_162.vcd");
  if(my_type==1 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_163.vcd");
  if(my_type==1 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_164.vcd");
  if(my_type==1 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_165.vcd");
  if(my_type==1 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_166.vcd");
  if(my_type==1 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_167.vcd");
  if(my_type==1 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_168.vcd");
  if(my_type==1 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_169.vcd");
  if(my_type==1 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_170.vcd");
  if(my_type==1 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_171.vcd");
  if(my_type==1 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_172.vcd");
  if(my_type==1 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_173.vcd");
  if(my_type==1 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_174.vcd");
  if(my_type==1 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_175.vcd");
  if(my_type==1 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_176.vcd");
  if(my_type==1 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_177.vcd");
  if(my_type==1 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_178.vcd");
  if(my_type==1 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_179.vcd");
  if(my_type==1 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_180.vcd");
  if(my_type==1 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_181.vcd");
  if(my_type==1 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_182.vcd");
  if(my_type==1 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_183.vcd");
  if(my_type==1 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_184.vcd");
  if(my_type==1 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_185.vcd");
  if(my_type==1 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_186.vcd");
  if(my_type==1 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_187.vcd");
  if(my_type==1 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_188.vcd");
  if(my_type==1 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_189.vcd");
  if(my_type==1 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_190.vcd");
  if(my_type==1 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_191.vcd");
  if(my_type==1 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_192.vcd");
  if(my_type==1 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_193.vcd");
  if(my_type==1 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_194.vcd");
  if(my_type==1 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_195.vcd");
  if(my_type==1 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_196.vcd");
  if(my_type==1 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_197.vcd");
  if(my_type==1 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_198.vcd");
  if(my_type==1 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_199.vcd");
  if(my_type==1 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_200.vcd");
  if(my_type==1 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_201.vcd");
  if(my_type==1 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_202.vcd");
  if(my_type==1 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_203.vcd");
  if(my_type==1 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_204.vcd");
  if(my_type==1 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_205.vcd");
  if(my_type==1 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_206.vcd");
  if(my_type==1 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_207.vcd");
  if(my_type==1 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_208.vcd");
  if(my_type==1 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_209.vcd");
  if(my_type==1 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_210.vcd");
  if(my_type==1 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_211.vcd");
  if(my_type==1 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_212.vcd");
  if(my_type==1 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_213.vcd");
  if(my_type==1 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_214.vcd");
  if(my_type==1 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_215.vcd");
  if(my_type==1 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_216.vcd");
  if(my_type==1 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_217.vcd");
  if(my_type==1 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_218.vcd");
  if(my_type==1 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_219.vcd");
  if(my_type==1 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_220.vcd");
  if(my_type==1 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_221.vcd");
  if(my_type==1 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_222.vcd");
  if(my_type==1 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_223.vcd");
  if(my_type==1 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_224.vcd");
  if(my_type==1 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_225.vcd");
  if(my_type==1 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_226.vcd");
  if(my_type==1 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_227.vcd");
  if(my_type==1 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_228.vcd");
  if(my_type==1 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_229.vcd");
  if(my_type==1 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_230.vcd");
  if(my_type==1 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_231.vcd");
  if(my_type==1 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_232.vcd");
  if(my_type==1 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_233.vcd");
  if(my_type==1 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_234.vcd");
  if(my_type==1 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_235.vcd");
  if(my_type==1 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_236.vcd");
  if(my_type==1 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_237.vcd");
  if(my_type==1 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_238.vcd");
  if(my_type==1 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_239.vcd");
  if(my_type==1 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_240.vcd");
  if(my_type==1 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_241.vcd");
  if(my_type==1 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_242.vcd");
  if(my_type==1 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_243.vcd");
  if(my_type==1 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_244.vcd");
  if(my_type==1 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_245.vcd");
  if(my_type==1 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_246.vcd");
  if(my_type==1 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_247.vcd");
  if(my_type==1 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_248.vcd");
  if(my_type==1 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_249.vcd");
  if(my_type==1 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_250.vcd");
  if(my_type==1 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_251.vcd");
  if(my_type==1 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_252.vcd");
  if(my_type==1 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_253.vcd");
  if(my_type==1 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_254.vcd");
  if(my_type==1 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_255.vcd");
  if(my_type==1 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_256.vcd");
  if(my_type==1 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_257.vcd");
  if(my_type==1 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_258.vcd");
  if(my_type==1 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_259.vcd");
  if(my_type==1 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_260.vcd");
  if(my_type==1 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_261.vcd");
  if(my_type==1 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_262.vcd");
  if(my_type==1 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_263.vcd");
  if(my_type==1 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_264.vcd");
  if(my_type==1 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_265.vcd");
  if(my_type==1 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_266.vcd");
  if(my_type==1 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_267.vcd");
  if(my_type==1 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_268.vcd");
  if(my_type==1 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_269.vcd");
  if(my_type==1 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_270.vcd");
  if(my_type==1 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_271.vcd");
  if(my_type==1 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_272.vcd");
  if(my_type==1 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_273.vcd");
  if(my_type==1 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_274.vcd");
  if(my_type==1 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_275.vcd");
  if(my_type==1 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_276.vcd");
  if(my_type==1 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_277.vcd");
  if(my_type==1 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_278.vcd");
  if(my_type==1 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_279.vcd");
  if(my_type==1 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_280.vcd");
  if(my_type==1 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_281.vcd");
  if(my_type==1 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_282.vcd");
  if(my_type==1 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_283.vcd");
  if(my_type==1 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_284.vcd");
  if(my_type==1 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_285.vcd");
  if(my_type==1 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_286.vcd");
  if(my_type==1 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_287.vcd");
  if(my_type==1 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_288.vcd");
  if(my_type==1 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_289.vcd");
  if(my_type==1 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_290.vcd");
  if(my_type==1 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_291.vcd");
  if(my_type==1 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_292.vcd");
  if(my_type==1 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_293.vcd");
  if(my_type==1 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_294.vcd");
  if(my_type==1 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_295.vcd");
  if(my_type==1 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_296.vcd");
  if(my_type==1 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_297.vcd");
  if(my_type==1 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_298.vcd");
  if(my_type==1 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_299.vcd");
  if(my_type==1 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_300.vcd");
  if(my_type==1 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_301.vcd");
  if(my_type==1 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_302.vcd");
  if(my_type==1 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_303.vcd");
  if(my_type==1 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_304.vcd");
  if(my_type==1 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_305.vcd");
  if(my_type==1 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_306.vcd");
  if(my_type==1 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_307.vcd");
  if(my_type==1 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_308.vcd");
  if(my_type==1 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_309.vcd");
  if(my_type==1 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_310.vcd");
  if(my_type==1 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_311.vcd");
  if(my_type==1 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_312.vcd");
  if(my_type==1 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_313.vcd");
  if(my_type==1 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_314.vcd");
  if(my_type==1 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_315.vcd");
  if(my_type==1 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_316.vcd");
  if(my_type==1 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_317.vcd");
  if(my_type==1 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_318.vcd");
  if(my_type==1 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_319.vcd");
  if(my_type==1 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_320.vcd");
  if(my_type==1 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_321.vcd");
  if(my_type==1 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_322.vcd");
  if(my_type==1 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_323.vcd");
  if(my_type==1 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_324.vcd");
  if(my_type==1 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_325.vcd");
  if(my_type==1 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_326.vcd");
  if(my_type==1 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_327.vcd");
  if(my_type==1 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_328.vcd");
  if(my_type==1 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_329.vcd");
  if(my_type==1 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_330.vcd");
  if(my_type==1 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_331.vcd");
  if(my_type==1 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_332.vcd");
  if(my_type==1 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_333.vcd");
  if(my_type==1 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_334.vcd");
  if(my_type==1 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_335.vcd");
  if(my_type==1 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_336.vcd");
  if(my_type==1 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_337.vcd");
  if(my_type==1 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_338.vcd");
  if(my_type==1 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_339.vcd");
  if(my_type==1 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_340.vcd");
  if(my_type==1 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_341.vcd");
  if(my_type==1 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_342.vcd");
  if(my_type==1 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_343.vcd");
  if(my_type==1 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_344.vcd");
  if(my_type==1 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_345.vcd");
  if(my_type==1 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_346.vcd");
  if(my_type==1 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_347.vcd");
  if(my_type==1 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_348.vcd");
  if(my_type==1 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_349.vcd");
  if(my_type==1 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_350.vcd");
  if(my_type==1 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_351.vcd");
  if(my_type==1 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_352.vcd");
  if(my_type==1 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_353.vcd");
  if(my_type==1 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_354.vcd");
  if(my_type==1 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_355.vcd");
  if(my_type==1 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_356.vcd");
  if(my_type==1 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_357.vcd");
  if(my_type==1 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_358.vcd");
  if(my_type==1 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_359.vcd");
  if(my_type==1 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_360.vcd");
  if(my_type==1 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_361.vcd");
  if(my_type==1 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_362.vcd");
  if(my_type==1 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_363.vcd");
  if(my_type==1 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_364.vcd");
  if(my_type==1 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_365.vcd");
  if(my_type==1 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_366.vcd");
  if(my_type==1 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_367.vcd");
  if(my_type==1 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_368.vcd");
  if(my_type==1 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_369.vcd");
  if(my_type==1 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_370.vcd");
  if(my_type==1 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_371.vcd");
  if(my_type==1 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_372.vcd");
  if(my_type==1 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_373.vcd");
  if(my_type==1 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_374.vcd");
  if(my_type==1 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_375.vcd");
  if(my_type==1 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_376.vcd");
  if(my_type==1 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_377.vcd");
  if(my_type==1 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_378.vcd");
  if(my_type==1 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_379.vcd");
  if(my_type==1 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_380.vcd");
  if(my_type==1 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_381.vcd");
  if(my_type==1 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_382.vcd");
  if(my_type==1 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_383.vcd");
  if(my_type==1 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_384.vcd");
  if(my_type==1 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_385.vcd");
  if(my_type==1 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_386.vcd");
  if(my_type==1 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_387.vcd");
  if(my_type==1 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_388.vcd");
  if(my_type==1 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_389.vcd");
  if(my_type==1 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_390.vcd");
  if(my_type==1 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_391.vcd");
  if(my_type==1 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_392.vcd");
  if(my_type==1 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_393.vcd");
  if(my_type==1 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_394.vcd");
  if(my_type==1 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_395.vcd");
  if(my_type==1 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_396.vcd");
  if(my_type==1 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_397.vcd");
  if(my_type==1 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_398.vcd");
  if(my_type==1 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_399.vcd");
  if(my_type==1 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_400.vcd");
  if(my_type==1 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_401.vcd");
  if(my_type==1 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_402.vcd");
  if(my_type==1 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_403.vcd");
  if(my_type==1 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_404.vcd");
  if(my_type==1 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_405.vcd");
  if(my_type==1 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_406.vcd");
  if(my_type==1 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_407.vcd");
  if(my_type==1 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_408.vcd");
  if(my_type==1 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_409.vcd");
  if(my_type==1 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_410.vcd");
  if(my_type==1 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_411.vcd");
  if(my_type==1 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_412.vcd");
  if(my_type==1 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_413.vcd");
  if(my_type==1 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_414.vcd");
  if(my_type==1 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_415.vcd");
  if(my_type==1 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_416.vcd");
  if(my_type==1 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_417.vcd");
  if(my_type==1 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_418.vcd");
  if(my_type==1 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_419.vcd");
  if(my_type==1 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_420.vcd");
  if(my_type==1 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_421.vcd");
  if(my_type==1 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_422.vcd");
  if(my_type==1 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_423.vcd");
  if(my_type==1 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_424.vcd");
  if(my_type==1 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_425.vcd");
  if(my_type==1 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_426.vcd");
  if(my_type==1 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_427.vcd");
  if(my_type==1 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_428.vcd");
  if(my_type==1 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_429.vcd");
  if(my_type==1 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_430.vcd");
  if(my_type==1 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_431.vcd");
  if(my_type==1 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_432.vcd");
  if(my_type==1 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_433.vcd");
  if(my_type==1 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_434.vcd");
  if(my_type==1 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_435.vcd");
  if(my_type==1 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_436.vcd");
  if(my_type==1 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_437.vcd");
  if(my_type==1 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_438.vcd");
  if(my_type==1 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_439.vcd");
  if(my_type==1 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_440.vcd");
  if(my_type==1 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_441.vcd");
  if(my_type==1 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_442.vcd");
  if(my_type==1 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_443.vcd");
  if(my_type==1 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_444.vcd");
  if(my_type==1 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_445.vcd");
  if(my_type==1 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_446.vcd");
  if(my_type==1 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_447.vcd");
  if(my_type==1 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_448.vcd");
  if(my_type==1 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_449.vcd");
  if(my_type==1 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_450.vcd");
  if(my_type==1 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_451.vcd");
  if(my_type==1 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_452.vcd");
  if(my_type==1 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_453.vcd");
  if(my_type==1 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_454.vcd");
  if(my_type==1 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_455.vcd");
  if(my_type==1 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_456.vcd");
  if(my_type==1 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_457.vcd");
  if(my_type==1 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_458.vcd");
  if(my_type==1 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_459.vcd");
  if(my_type==1 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_460.vcd");
  if(my_type==1 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_461.vcd");
  if(my_type==1 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_462.vcd");
  if(my_type==1 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_463.vcd");
  if(my_type==1 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_464.vcd");
  if(my_type==1 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_465.vcd");
  if(my_type==1 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_466.vcd");
  if(my_type==1 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_467.vcd");
  if(my_type==1 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_468.vcd");
  if(my_type==1 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_469.vcd");
  if(my_type==1 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_470.vcd");
  if(my_type==1 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_471.vcd");
  if(my_type==1 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_472.vcd");
  if(my_type==1 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_473.vcd");
  if(my_type==1 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_474.vcd");
  if(my_type==1 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_475.vcd");
  if(my_type==1 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_476.vcd");
  if(my_type==1 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_477.vcd");
  if(my_type==1 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_478.vcd");
  if(my_type==1 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_479.vcd");
  if(my_type==1 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_480.vcd");
  if(my_type==1 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_481.vcd");
  if(my_type==1 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_482.vcd");
  if(my_type==1 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_483.vcd");
  if(my_type==1 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_484.vcd");
  if(my_type==1 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_485.vcd");
  if(my_type==1 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_486.vcd");
  if(my_type==1 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_487.vcd");
  if(my_type==1 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_488.vcd");
  if(my_type==1 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_489.vcd");
  if(my_type==1 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_490.vcd");
  if(my_type==1 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_491.vcd");
  if(my_type==1 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_492.vcd");
  if(my_type==1 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_493.vcd");
  if(my_type==1 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_494.vcd");
  if(my_type==1 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_495.vcd");
  if(my_type==1 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_496.vcd");
  if(my_type==1 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_497.vcd");
  if(my_type==1 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_498.vcd");
  if(my_type==1 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_499.vcd");
  if(my_type==1 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_500.vcd");
  if(my_type==1 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_501.vcd");
  if(my_type==1 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_502.vcd");
  if(my_type==1 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_503.vcd");
  if(my_type==1 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_504.vcd");
  if(my_type==1 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_505.vcd");
  if(my_type==1 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_506.vcd");
  if(my_type==1 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_507.vcd");
  if(my_type==1 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_508.vcd");
  if(my_type==1 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_509.vcd");
  if(my_type==1 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_510.vcd");
  if(my_type==1 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_511.vcd");
  if(my_type==1 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_512.vcd");
  if(my_type==1 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_513.vcd");
  if(my_type==1 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_514.vcd");
  if(my_type==1 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_515.vcd");
  if(my_type==1 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_516.vcd");
  if(my_type==1 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_517.vcd");
  if(my_type==1 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_518.vcd");
  if(my_type==1 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_519.vcd");
  if(my_type==1 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_520.vcd");
  if(my_type==1 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_521.vcd");
  if(my_type==1 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_522.vcd");
  if(my_type==1 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_523.vcd");
  if(my_type==1 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_524.vcd");
  if(my_type==1 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_525.vcd");
  if(my_type==1 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_526.vcd");
  if(my_type==1 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_527.vcd");
  if(my_type==1 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_528.vcd");
  if(my_type==1 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_529.vcd");
  if(my_type==1 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_530.vcd");
  if(my_type==1 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_531.vcd");
  if(my_type==1 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_532.vcd");
  if(my_type==1 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_533.vcd");
  if(my_type==1 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_534.vcd");
  if(my_type==1 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_535.vcd");
  if(my_type==1 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_536.vcd");
  if(my_type==1 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_537.vcd");
  if(my_type==1 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_538.vcd");
  if(my_type==1 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_539.vcd");
  if(my_type==1 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_540.vcd");
  if(my_type==1 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_541.vcd");
  if(my_type==1 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_542.vcd");
  if(my_type==1 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_543.vcd");
  if(my_type==1 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_544.vcd");
  if(my_type==1 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_545.vcd");
  if(my_type==1 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_546.vcd");
  if(my_type==1 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_547.vcd");
  if(my_type==1 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_548.vcd");
  if(my_type==1 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_549.vcd");
  if(my_type==1 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_550.vcd");
  if(my_type==1 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_551.vcd");
  if(my_type==1 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_552.vcd");
  if(my_type==1 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_553.vcd");
  if(my_type==1 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_554.vcd");
  if(my_type==1 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_555.vcd");
  if(my_type==1 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_556.vcd");
  if(my_type==1 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_557.vcd");
  if(my_type==1 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_558.vcd");
  if(my_type==1 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_559.vcd");
  if(my_type==1 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_560.vcd");
  if(my_type==1 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_561.vcd");
  if(my_type==1 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_562.vcd");
  if(my_type==1 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_563.vcd");
  if(my_type==1 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_564.vcd");
  if(my_type==1 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_565.vcd");
  if(my_type==1 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_566.vcd");
  if(my_type==1 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_567.vcd");
  if(my_type==1 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_568.vcd");
  if(my_type==1 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_569.vcd");
  if(my_type==1 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_570.vcd");
  if(my_type==1 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_571.vcd");
  if(my_type==1 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_572.vcd");
  if(my_type==1 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_573.vcd");
  if(my_type==1 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_574.vcd");
  if(my_type==1 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_575.vcd");
  if(my_type==1 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_576.vcd");
  if(my_type==1 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_577.vcd");
  if(my_type==1 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_578.vcd");
  if(my_type==1 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_579.vcd");
  if(my_type==1 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_580.vcd");
  if(my_type==1 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_581.vcd");
  if(my_type==1 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_582.vcd");
  if(my_type==1 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_583.vcd");
  if(my_type==1 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_584.vcd");
  if(my_type==1 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_585.vcd");
  if(my_type==1 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_586.vcd");
  if(my_type==1 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_587.vcd");
  if(my_type==1 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_588.vcd");
  if(my_type==1 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_589.vcd");
  if(my_type==1 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_590.vcd");
  if(my_type==1 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_591.vcd");
  if(my_type==1 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_592.vcd");
  if(my_type==1 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_593.vcd");
  if(my_type==1 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_594.vcd");
  if(my_type==1 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_595.vcd");
  if(my_type==1 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_596.vcd");
  if(my_type==1 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_597.vcd");
  if(my_type==1 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_598.vcd");
  if(my_type==1 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_599.vcd");
  if(my_type==1 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_600.vcd");
  if(my_type==1 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_601.vcd");
  if(my_type==1 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_602.vcd");
  if(my_type==1 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_603.vcd");
  if(my_type==1 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_604.vcd");
  if(my_type==1 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_605.vcd");
  if(my_type==1 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_606.vcd");
  if(my_type==1 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_607.vcd");
  if(my_type==1 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_608.vcd");
  if(my_type==1 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_609.vcd");
  if(my_type==1 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_610.vcd");
  if(my_type==1 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_611.vcd");
  if(my_type==1 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_612.vcd");
  if(my_type==1 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_613.vcd");
  if(my_type==1 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_614.vcd");
  if(my_type==1 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_615.vcd");
  if(my_type==1 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_616.vcd");
  if(my_type==1 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_617.vcd");
  if(my_type==1 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_618.vcd");
  if(my_type==1 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_619.vcd");
  if(my_type==1 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_620.vcd");
  if(my_type==1 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_621.vcd");
  if(my_type==1 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_622.vcd");
  if(my_type==1 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_623.vcd");
  if(my_type==1 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_624.vcd");
  if(my_type==1 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_625.vcd");
  if(my_type==1 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_626.vcd");
  if(my_type==1 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_627.vcd");
  if(my_type==1 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_628.vcd");
  if(my_type==1 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_629.vcd");
  if(my_type==1 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_630.vcd");
  if(my_type==1 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_631.vcd");
  if(my_type==1 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_632.vcd");
  if(my_type==1 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_633.vcd");
  if(my_type==1 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_634.vcd");
  if(my_type==1 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_635.vcd");
  if(my_type==1 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_636.vcd");
  if(my_type==1 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_637.vcd");
  if(my_type==1 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_638.vcd");
  if(my_type==1 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_639.vcd");
  if(my_type==1 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_640.vcd");
  if(my_type==1 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_641.vcd");
  if(my_type==1 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_642.vcd");
  if(my_type==1 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_643.vcd");
  if(my_type==1 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_644.vcd");
  if(my_type==1 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_645.vcd");
  if(my_type==1 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_646.vcd");
  if(my_type==1 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_647.vcd");
  if(my_type==1 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_648.vcd");
  if(my_type==1 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_649.vcd");
  if(my_type==1 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_650.vcd");
  if(my_type==1 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_651.vcd");
  if(my_type==1 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_652.vcd");
  if(my_type==1 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_653.vcd");
  if(my_type==1 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_654.vcd");
  if(my_type==1 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_655.vcd");
  if(my_type==1 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_656.vcd");
  if(my_type==1 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_657.vcd");
  if(my_type==1 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_658.vcd");
  if(my_type==1 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_659.vcd");
  if(my_type==1 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_660.vcd");
  if(my_type==1 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_661.vcd");
  if(my_type==1 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_662.vcd");
  if(my_type==1 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_663.vcd");
  if(my_type==1 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_664.vcd");
  if(my_type==1 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_665.vcd");
  if(my_type==1 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_666.vcd");
  if(my_type==1 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_667.vcd");
  if(my_type==1 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_668.vcd");
  if(my_type==1 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_669.vcd");
  if(my_type==1 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_670.vcd");
  if(my_type==1 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_671.vcd");
  if(my_type==1 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_672.vcd");
  if(my_type==1 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_673.vcd");
  if(my_type==1 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_674.vcd");
  if(my_type==1 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_675.vcd");
  if(my_type==1 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_676.vcd");
  if(my_type==1 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_677.vcd");
  if(my_type==1 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_678.vcd");
  if(my_type==1 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_679.vcd");
  if(my_type==1 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_680.vcd");
  if(my_type==1 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_681.vcd");
  if(my_type==1 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_682.vcd");
  if(my_type==1 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_683.vcd");
  if(my_type==1 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_684.vcd");
  if(my_type==1 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_685.vcd");
  if(my_type==1 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_686.vcd");
  if(my_type==1 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_687.vcd");
  if(my_type==1 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_688.vcd");
  if(my_type==1 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_689.vcd");
  if(my_type==1 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_690.vcd");
  if(my_type==1 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_691.vcd");
  if(my_type==1 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_692.vcd");
  if(my_type==1 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_693.vcd");
  if(my_type==1 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_694.vcd");
  if(my_type==1 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_695.vcd");
  if(my_type==1 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_696.vcd");
  if(my_type==1 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_697.vcd");
  if(my_type==1 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_698.vcd");
  if(my_type==1 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_699.vcd");
  if(my_type==1 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_700.vcd");
  if(my_type==1 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_701.vcd");
  if(my_type==1 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_702.vcd");
  if(my_type==1 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_703.vcd");
  if(my_type==1 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_704.vcd");
  if(my_type==1 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_705.vcd");
  if(my_type==1 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_706.vcd");
  if(my_type==1 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_707.vcd");
  if(my_type==1 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_708.vcd");
  if(my_type==1 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_709.vcd");
  if(my_type==1 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_710.vcd");
  if(my_type==1 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_711.vcd");
  if(my_type==1 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_712.vcd");
  if(my_type==1 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_713.vcd");
  if(my_type==1 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_714.vcd");
  if(my_type==1 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_715.vcd");
  if(my_type==1 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_716.vcd");
  if(my_type==1 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_717.vcd");
  if(my_type==1 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_718.vcd");
  if(my_type==1 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_719.vcd");
  if(my_type==1 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_720.vcd");
  if(my_type==1 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_721.vcd");
  if(my_type==1 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_722.vcd");
  if(my_type==1 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_723.vcd");
  if(my_type==1 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_724.vcd");
  if(my_type==1 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_725.vcd");
  if(my_type==1 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_726.vcd");
  if(my_type==1 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_727.vcd");
  if(my_type==1 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_728.vcd");
  if(my_type==1 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_729.vcd");
  if(my_type==1 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_730.vcd");
  if(my_type==1 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_731.vcd");
  if(my_type==1 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_732.vcd");
  if(my_type==1 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_733.vcd");
  if(my_type==1 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_734.vcd");
  if(my_type==1 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_735.vcd");
  if(my_type==1 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_736.vcd");
  if(my_type==1 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_737.vcd");
  if(my_type==1 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_738.vcd");
  if(my_type==1 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_739.vcd");
  if(my_type==1 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_740.vcd");
  if(my_type==1 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_741.vcd");
  if(my_type==1 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_742.vcd");
  if(my_type==1 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_743.vcd");
  if(my_type==1 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_744.vcd");
  if(my_type==1 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_745.vcd");
  if(my_type==1 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_746.vcd");
  if(my_type==1 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_747.vcd");
  if(my_type==1 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_748.vcd");
  if(my_type==1 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_749.vcd");
  if(my_type==1 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_750.vcd");
  if(my_type==1 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_751.vcd");
  if(my_type==1 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_752.vcd");
  if(my_type==1 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_753.vcd");
  if(my_type==1 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_754.vcd");
  if(my_type==1 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_755.vcd");
  if(my_type==1 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_756.vcd");
  if(my_type==1 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_757.vcd");
  if(my_type==1 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_758.vcd");
  if(my_type==1 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_759.vcd");
  if(my_type==1 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_760.vcd");
  if(my_type==1 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_761.vcd");
  if(my_type==1 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_762.vcd");
  if(my_type==1 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_763.vcd");
  if(my_type==1 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_764.vcd");
  if(my_type==1 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_765.vcd");
  if(my_type==1 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_766.vcd");
  if(my_type==1 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_767.vcd");
  if(my_type==1 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_768.vcd");
  if(my_type==1 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_769.vcd");
  if(my_type==1 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_770.vcd");
  if(my_type==1 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_771.vcd");
  if(my_type==1 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_772.vcd");
  if(my_type==1 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_773.vcd");
  if(my_type==1 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_774.vcd");
  if(my_type==1 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_775.vcd");
  if(my_type==1 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_776.vcd");
  if(my_type==1 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_777.vcd");
  if(my_type==1 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_778.vcd");
  if(my_type==1 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_779.vcd");
  if(my_type==1 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_780.vcd");
  if(my_type==1 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_781.vcd");
  if(my_type==1 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_782.vcd");
  if(my_type==1 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_783.vcd");
  if(my_type==1 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_784.vcd");
  if(my_type==1 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_785.vcd");
  if(my_type==1 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_786.vcd");
  if(my_type==1 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_787.vcd");
  if(my_type==1 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_788.vcd");
  if(my_type==1 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_789.vcd");
  if(my_type==1 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_790.vcd");
  if(my_type==1 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_791.vcd");
  if(my_type==1 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_792.vcd");
  if(my_type==1 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_793.vcd");
  if(my_type==1 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_794.vcd");
  if(my_type==1 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_795.vcd");
  if(my_type==1 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_796.vcd");
  if(my_type==1 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_797.vcd");
  if(my_type==1 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_798.vcd");
  if(my_type==1 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_799.vcd");
  if(my_type==1 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_800.vcd");
  if(my_type==1 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_801.vcd");
  if(my_type==1 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_802.vcd");
  if(my_type==1 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_803.vcd");
  if(my_type==1 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_804.vcd");
  if(my_type==1 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_805.vcd");
  if(my_type==1 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_806.vcd");
  if(my_type==1 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_807.vcd");
  if(my_type==1 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_808.vcd");
  if(my_type==1 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_809.vcd");
  if(my_type==1 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_810.vcd");
  if(my_type==1 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_811.vcd");
  if(my_type==1 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_812.vcd");
  if(my_type==1 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_813.vcd");
  if(my_type==1 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_814.vcd");
  if(my_type==1 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_815.vcd");
  if(my_type==1 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_816.vcd");
  if(my_type==1 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_817.vcd");
  if(my_type==1 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_818.vcd");
  if(my_type==1 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_819.vcd");
  if(my_type==1 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_820.vcd");
  if(my_type==1 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_821.vcd");
  if(my_type==1 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_822.vcd");
  if(my_type==1 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_823.vcd");
  if(my_type==1 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_824.vcd");
  if(my_type==1 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_825.vcd");
  if(my_type==1 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_826.vcd");
  if(my_type==1 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_827.vcd");
  if(my_type==1 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_828.vcd");
  if(my_type==1 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_829.vcd");
  if(my_type==1 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_830.vcd");
  if(my_type==1 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_831.vcd");
  if(my_type==1 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_832.vcd");
  if(my_type==1 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_833.vcd");
  if(my_type==1 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_834.vcd");
  if(my_type==1 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_835.vcd");
  if(my_type==1 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_836.vcd");
  if(my_type==1 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_837.vcd");
  if(my_type==1 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_838.vcd");
  if(my_type==1 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_839.vcd");
  if(my_type==1 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_840.vcd");
  if(my_type==1 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_841.vcd");
  if(my_type==1 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_842.vcd");
  if(my_type==1 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_843.vcd");
  if(my_type==1 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_844.vcd");
  if(my_type==1 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_845.vcd");
  if(my_type==1 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_846.vcd");
  if(my_type==1 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_847.vcd");
  if(my_type==1 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_848.vcd");
  if(my_type==1 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_849.vcd");
  if(my_type==1 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_850.vcd");
  if(my_type==1 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_851.vcd");
  if(my_type==1 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_852.vcd");
  if(my_type==1 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_853.vcd");
  if(my_type==1 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_854.vcd");
  if(my_type==1 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_855.vcd");
  if(my_type==1 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_856.vcd");
  if(my_type==1 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_857.vcd");
  if(my_type==1 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_858.vcd");
  if(my_type==1 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_859.vcd");
  if(my_type==1 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_860.vcd");
  if(my_type==1 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_861.vcd");
  if(my_type==1 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_862.vcd");
  if(my_type==1 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_863.vcd");
  if(my_type==1 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_864.vcd");
  if(my_type==1 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_865.vcd");
  if(my_type==1 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_866.vcd");
  if(my_type==1 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_867.vcd");
  if(my_type==1 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_868.vcd");
  if(my_type==1 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_869.vcd");
  if(my_type==1 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_870.vcd");
  if(my_type==1 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_871.vcd");
  if(my_type==1 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_872.vcd");
  if(my_type==1 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_873.vcd");
  if(my_type==1 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_874.vcd");
  if(my_type==1 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_875.vcd");
  if(my_type==1 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_876.vcd");
  if(my_type==1 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_877.vcd");
  if(my_type==1 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_878.vcd");
  if(my_type==1 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_879.vcd");
  if(my_type==1 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_880.vcd");
  if(my_type==1 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_881.vcd");
  if(my_type==1 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_882.vcd");
  if(my_type==1 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_883.vcd");
  if(my_type==1 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_884.vcd");
  if(my_type==1 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_885.vcd");
  if(my_type==1 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_886.vcd");
  if(my_type==1 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_887.vcd");
  if(my_type==1 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_888.vcd");
  if(my_type==1 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_889.vcd");
  if(my_type==1 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_890.vcd");
  if(my_type==1 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_891.vcd");
  if(my_type==1 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_892.vcd");
  if(my_type==1 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_893.vcd");
  if(my_type==1 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_894.vcd");
  if(my_type==1 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_895.vcd");
  if(my_type==1 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_896.vcd");
  if(my_type==1 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_897.vcd");
  if(my_type==1 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_898.vcd");
  if(my_type==1 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_899.vcd");
  if(my_type==1 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_900.vcd");
  if(my_type==1 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_901.vcd");
  if(my_type==1 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_902.vcd");
  if(my_type==1 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_903.vcd");
  if(my_type==1 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_904.vcd");
  if(my_type==1 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_905.vcd");
  if(my_type==1 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_906.vcd");
  if(my_type==1 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_907.vcd");
  if(my_type==1 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_908.vcd");
  if(my_type==1 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_909.vcd");
  if(my_type==1 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_910.vcd");
  if(my_type==1 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_911.vcd");
  if(my_type==1 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_912.vcd");
  if(my_type==1 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_913.vcd");
  if(my_type==1 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_914.vcd");
  if(my_type==1 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_915.vcd");
  if(my_type==1 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_916.vcd");
  if(my_type==1 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_917.vcd");
  if(my_type==1 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_918.vcd");
  if(my_type==1 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_919.vcd");
  if(my_type==1 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_920.vcd");
  if(my_type==1 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_921.vcd");
  if(my_type==1 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_922.vcd");
  if(my_type==1 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_923.vcd");
  if(my_type==1 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_924.vcd");
  if(my_type==1 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_925.vcd");
  if(my_type==1 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_926.vcd");
  if(my_type==1 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_927.vcd");
  if(my_type==1 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_928.vcd");
  if(my_type==1 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_929.vcd");
  if(my_type==1 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_930.vcd");
  if(my_type==1 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_931.vcd");
  if(my_type==1 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_932.vcd");
  if(my_type==1 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_933.vcd");
  if(my_type==1 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_934.vcd");
  if(my_type==1 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_935.vcd");
  if(my_type==1 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_936.vcd");
  if(my_type==1 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_937.vcd");
  if(my_type==1 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_938.vcd");
  if(my_type==1 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_939.vcd");
  if(my_type==1 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_940.vcd");
  if(my_type==1 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_941.vcd");
  if(my_type==1 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_942.vcd");
  if(my_type==1 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_943.vcd");
  if(my_type==1 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_944.vcd");
  if(my_type==1 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_945.vcd");
  if(my_type==1 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_946.vcd");
  if(my_type==1 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_947.vcd");
  if(my_type==1 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_948.vcd");
  if(my_type==1 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_949.vcd");
  if(my_type==1 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_950.vcd");
  if(my_type==1 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_951.vcd");
  if(my_type==1 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_952.vcd");
  if(my_type==1 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_953.vcd");
  if(my_type==1 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_954.vcd");
  if(my_type==1 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_955.vcd");
  if(my_type==1 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_956.vcd");
  if(my_type==1 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_957.vcd");
  if(my_type==1 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_958.vcd");
  if(my_type==1 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_959.vcd");
  if(my_type==1 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_960.vcd");
  if(my_type==1 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_961.vcd");
  if(my_type==1 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_962.vcd");
  if(my_type==1 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_963.vcd");
  if(my_type==1 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_964.vcd");
  if(my_type==1 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_965.vcd");
  if(my_type==1 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_966.vcd");
  if(my_type==1 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_967.vcd");
  if(my_type==1 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_968.vcd");
  if(my_type==1 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_969.vcd");
  if(my_type==1 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_970.vcd");
  if(my_type==1 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_971.vcd");
  if(my_type==1 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_972.vcd");
  if(my_type==1 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_973.vcd");
  if(my_type==1 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_974.vcd");
  if(my_type==1 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_975.vcd");
  if(my_type==1 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_976.vcd");
  if(my_type==1 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_977.vcd");
  if(my_type==1 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_978.vcd");
  if(my_type==1 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_979.vcd");
  if(my_type==1 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_980.vcd");
  if(my_type==1 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_981.vcd");
  if(my_type==1 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_982.vcd");
  if(my_type==1 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_983.vcd");
  if(my_type==1 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_984.vcd");
  if(my_type==1 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_985.vcd");
  if(my_type==1 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_986.vcd");
  if(my_type==1 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_987.vcd");
  if(my_type==1 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_988.vcd");
  if(my_type==1 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_989.vcd");
  if(my_type==1 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_990.vcd");
  if(my_type==1 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_991.vcd");
  if(my_type==1 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_992.vcd");
  if(my_type==1 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_993.vcd");
  if(my_type==1 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_994.vcd");
  if(my_type==1 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_995.vcd");
  if(my_type==1 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_996.vcd");
  if(my_type==1 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_997.vcd");
  if(my_type==1 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_998.vcd");
  if(my_type==1 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_1_999.vcd");
  if(my_type==2 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_0.vcd");
  if(my_type==2 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_1.vcd");
  if(my_type==2 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_2.vcd");
  if(my_type==2 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_3.vcd");
  if(my_type==2 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_4.vcd");
  if(my_type==2 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_5.vcd");
  if(my_type==2 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_6.vcd");
  if(my_type==2 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_7.vcd");
  if(my_type==2 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_8.vcd");
  if(my_type==2 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_9.vcd");
  if(my_type==2 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_10.vcd");
  if(my_type==2 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_11.vcd");
  if(my_type==2 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_12.vcd");
  if(my_type==2 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_13.vcd");
  if(my_type==2 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_14.vcd");
  if(my_type==2 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_15.vcd");
  if(my_type==2 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_16.vcd");
  if(my_type==2 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_17.vcd");
  if(my_type==2 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_18.vcd");
  if(my_type==2 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_19.vcd");
  if(my_type==2 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_20.vcd");
  if(my_type==2 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_21.vcd");
  if(my_type==2 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_22.vcd");
  if(my_type==2 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_23.vcd");
  if(my_type==2 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_24.vcd");
  if(my_type==2 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_25.vcd");
  if(my_type==2 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_26.vcd");
  if(my_type==2 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_27.vcd");
  if(my_type==2 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_28.vcd");
  if(my_type==2 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_29.vcd");
  if(my_type==2 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_30.vcd");
  if(my_type==2 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_31.vcd");
  if(my_type==2 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_32.vcd");
  if(my_type==2 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_33.vcd");
  if(my_type==2 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_34.vcd");
  if(my_type==2 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_35.vcd");
  if(my_type==2 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_36.vcd");
  if(my_type==2 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_37.vcd");
  if(my_type==2 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_38.vcd");
  if(my_type==2 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_39.vcd");
  if(my_type==2 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_40.vcd");
  if(my_type==2 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_41.vcd");
  if(my_type==2 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_42.vcd");
  if(my_type==2 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_43.vcd");
  if(my_type==2 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_44.vcd");
  if(my_type==2 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_45.vcd");
  if(my_type==2 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_46.vcd");
  if(my_type==2 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_47.vcd");
  if(my_type==2 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_48.vcd");
  if(my_type==2 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_49.vcd");
  if(my_type==2 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_50.vcd");
  if(my_type==2 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_51.vcd");
  if(my_type==2 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_52.vcd");
  if(my_type==2 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_53.vcd");
  if(my_type==2 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_54.vcd");
  if(my_type==2 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_55.vcd");
  if(my_type==2 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_56.vcd");
  if(my_type==2 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_57.vcd");
  if(my_type==2 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_58.vcd");
  if(my_type==2 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_59.vcd");
  if(my_type==2 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_60.vcd");
  if(my_type==2 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_61.vcd");
  if(my_type==2 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_62.vcd");
  if(my_type==2 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_63.vcd");
  if(my_type==2 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_64.vcd");
  if(my_type==2 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_65.vcd");
  if(my_type==2 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_66.vcd");
  if(my_type==2 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_67.vcd");
  if(my_type==2 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_68.vcd");
  if(my_type==2 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_69.vcd");
  if(my_type==2 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_70.vcd");
  if(my_type==2 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_71.vcd");
  if(my_type==2 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_72.vcd");
  if(my_type==2 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_73.vcd");
  if(my_type==2 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_74.vcd");
  if(my_type==2 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_75.vcd");
  if(my_type==2 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_76.vcd");
  if(my_type==2 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_77.vcd");
  if(my_type==2 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_78.vcd");
  if(my_type==2 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_79.vcd");
  if(my_type==2 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_80.vcd");
  if(my_type==2 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_81.vcd");
  if(my_type==2 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_82.vcd");
  if(my_type==2 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_83.vcd");
  if(my_type==2 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_84.vcd");
  if(my_type==2 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_85.vcd");
  if(my_type==2 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_86.vcd");
  if(my_type==2 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_87.vcd");
  if(my_type==2 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_88.vcd");
  if(my_type==2 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_89.vcd");
  if(my_type==2 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_90.vcd");
  if(my_type==2 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_91.vcd");
  if(my_type==2 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_92.vcd");
  if(my_type==2 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_93.vcd");
  if(my_type==2 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_94.vcd");
  if(my_type==2 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_95.vcd");
  if(my_type==2 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_96.vcd");
  if(my_type==2 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_97.vcd");
  if(my_type==2 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_98.vcd");
  if(my_type==2 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_99.vcd");
  if(my_type==2 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_100.vcd");
  if(my_type==2 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_101.vcd");
  if(my_type==2 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_102.vcd");
  if(my_type==2 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_103.vcd");
  if(my_type==2 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_104.vcd");
  if(my_type==2 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_105.vcd");
  if(my_type==2 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_106.vcd");
  if(my_type==2 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_107.vcd");
  if(my_type==2 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_108.vcd");
  if(my_type==2 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_109.vcd");
  if(my_type==2 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_110.vcd");
  if(my_type==2 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_111.vcd");
  if(my_type==2 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_112.vcd");
  if(my_type==2 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_113.vcd");
  if(my_type==2 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_114.vcd");
  if(my_type==2 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_115.vcd");
  if(my_type==2 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_116.vcd");
  if(my_type==2 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_117.vcd");
  if(my_type==2 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_118.vcd");
  if(my_type==2 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_119.vcd");
  if(my_type==2 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_120.vcd");
  if(my_type==2 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_121.vcd");
  if(my_type==2 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_122.vcd");
  if(my_type==2 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_123.vcd");
  if(my_type==2 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_124.vcd");
  if(my_type==2 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_125.vcd");
  if(my_type==2 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_126.vcd");
  if(my_type==2 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_127.vcd");
  if(my_type==2 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_128.vcd");
  if(my_type==2 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_129.vcd");
  if(my_type==2 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_130.vcd");
  if(my_type==2 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_131.vcd");
  if(my_type==2 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_132.vcd");
  if(my_type==2 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_133.vcd");
  if(my_type==2 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_134.vcd");
  if(my_type==2 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_135.vcd");
  if(my_type==2 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_136.vcd");
  if(my_type==2 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_137.vcd");
  if(my_type==2 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_138.vcd");
  if(my_type==2 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_139.vcd");
  if(my_type==2 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_140.vcd");
  if(my_type==2 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_141.vcd");
  if(my_type==2 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_142.vcd");
  if(my_type==2 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_143.vcd");
  if(my_type==2 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_144.vcd");
  if(my_type==2 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_145.vcd");
  if(my_type==2 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_146.vcd");
  if(my_type==2 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_147.vcd");
  if(my_type==2 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_148.vcd");
  if(my_type==2 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_149.vcd");
  if(my_type==2 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_150.vcd");
  if(my_type==2 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_151.vcd");
  if(my_type==2 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_152.vcd");
  if(my_type==2 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_153.vcd");
  if(my_type==2 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_154.vcd");
  if(my_type==2 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_155.vcd");
  if(my_type==2 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_156.vcd");
  if(my_type==2 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_157.vcd");
  if(my_type==2 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_158.vcd");
  if(my_type==2 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_159.vcd");
  if(my_type==2 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_160.vcd");
  if(my_type==2 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_161.vcd");
  if(my_type==2 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_162.vcd");
  if(my_type==2 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_163.vcd");
  if(my_type==2 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_164.vcd");
  if(my_type==2 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_165.vcd");
  if(my_type==2 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_166.vcd");
  if(my_type==2 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_167.vcd");
  if(my_type==2 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_168.vcd");
  if(my_type==2 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_169.vcd");
  if(my_type==2 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_170.vcd");
  if(my_type==2 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_171.vcd");
  if(my_type==2 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_172.vcd");
  if(my_type==2 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_173.vcd");
  if(my_type==2 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_174.vcd");
  if(my_type==2 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_175.vcd");
  if(my_type==2 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_176.vcd");
  if(my_type==2 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_177.vcd");
  if(my_type==2 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_178.vcd");
  if(my_type==2 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_179.vcd");
  if(my_type==2 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_180.vcd");
  if(my_type==2 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_181.vcd");
  if(my_type==2 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_182.vcd");
  if(my_type==2 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_183.vcd");
  if(my_type==2 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_184.vcd");
  if(my_type==2 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_185.vcd");
  if(my_type==2 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_186.vcd");
  if(my_type==2 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_187.vcd");
  if(my_type==2 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_188.vcd");
  if(my_type==2 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_189.vcd");
  if(my_type==2 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_190.vcd");
  if(my_type==2 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_191.vcd");
  if(my_type==2 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_192.vcd");
  if(my_type==2 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_193.vcd");
  if(my_type==2 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_194.vcd");
  if(my_type==2 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_195.vcd");
  if(my_type==2 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_196.vcd");
  if(my_type==2 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_197.vcd");
  if(my_type==2 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_198.vcd");
  if(my_type==2 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_199.vcd");
  if(my_type==2 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_200.vcd");
  if(my_type==2 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_201.vcd");
  if(my_type==2 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_202.vcd");
  if(my_type==2 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_203.vcd");
  if(my_type==2 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_204.vcd");
  if(my_type==2 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_205.vcd");
  if(my_type==2 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_206.vcd");
  if(my_type==2 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_207.vcd");
  if(my_type==2 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_208.vcd");
  if(my_type==2 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_209.vcd");
  if(my_type==2 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_210.vcd");
  if(my_type==2 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_211.vcd");
  if(my_type==2 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_212.vcd");
  if(my_type==2 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_213.vcd");
  if(my_type==2 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_214.vcd");
  if(my_type==2 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_215.vcd");
  if(my_type==2 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_216.vcd");
  if(my_type==2 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_217.vcd");
  if(my_type==2 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_218.vcd");
  if(my_type==2 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_219.vcd");
  if(my_type==2 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_220.vcd");
  if(my_type==2 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_221.vcd");
  if(my_type==2 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_222.vcd");
  if(my_type==2 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_223.vcd");
  if(my_type==2 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_224.vcd");
  if(my_type==2 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_225.vcd");
  if(my_type==2 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_226.vcd");
  if(my_type==2 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_227.vcd");
  if(my_type==2 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_228.vcd");
  if(my_type==2 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_229.vcd");
  if(my_type==2 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_230.vcd");
  if(my_type==2 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_231.vcd");
  if(my_type==2 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_232.vcd");
  if(my_type==2 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_233.vcd");
  if(my_type==2 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_234.vcd");
  if(my_type==2 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_235.vcd");
  if(my_type==2 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_236.vcd");
  if(my_type==2 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_237.vcd");
  if(my_type==2 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_238.vcd");
  if(my_type==2 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_239.vcd");
  if(my_type==2 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_240.vcd");
  if(my_type==2 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_241.vcd");
  if(my_type==2 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_242.vcd");
  if(my_type==2 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_243.vcd");
  if(my_type==2 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_244.vcd");
  if(my_type==2 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_245.vcd");
  if(my_type==2 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_246.vcd");
  if(my_type==2 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_247.vcd");
  if(my_type==2 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_248.vcd");
  if(my_type==2 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_249.vcd");
  if(my_type==2 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_250.vcd");
  if(my_type==2 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_251.vcd");
  if(my_type==2 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_252.vcd");
  if(my_type==2 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_253.vcd");
  if(my_type==2 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_254.vcd");
  if(my_type==2 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_255.vcd");
  if(my_type==2 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_256.vcd");
  if(my_type==2 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_257.vcd");
  if(my_type==2 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_258.vcd");
  if(my_type==2 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_259.vcd");
  if(my_type==2 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_260.vcd");
  if(my_type==2 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_261.vcd");
  if(my_type==2 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_262.vcd");
  if(my_type==2 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_263.vcd");
  if(my_type==2 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_264.vcd");
  if(my_type==2 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_265.vcd");
  if(my_type==2 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_266.vcd");
  if(my_type==2 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_267.vcd");
  if(my_type==2 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_268.vcd");
  if(my_type==2 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_269.vcd");
  if(my_type==2 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_270.vcd");
  if(my_type==2 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_271.vcd");
  if(my_type==2 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_272.vcd");
  if(my_type==2 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_273.vcd");
  if(my_type==2 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_274.vcd");
  if(my_type==2 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_275.vcd");
  if(my_type==2 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_276.vcd");
  if(my_type==2 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_277.vcd");
  if(my_type==2 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_278.vcd");
  if(my_type==2 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_279.vcd");
  if(my_type==2 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_280.vcd");
  if(my_type==2 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_281.vcd");
  if(my_type==2 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_282.vcd");
  if(my_type==2 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_283.vcd");
  if(my_type==2 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_284.vcd");
  if(my_type==2 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_285.vcd");
  if(my_type==2 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_286.vcd");
  if(my_type==2 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_287.vcd");
  if(my_type==2 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_288.vcd");
  if(my_type==2 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_289.vcd");
  if(my_type==2 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_290.vcd");
  if(my_type==2 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_291.vcd");
  if(my_type==2 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_292.vcd");
  if(my_type==2 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_293.vcd");
  if(my_type==2 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_294.vcd");
  if(my_type==2 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_295.vcd");
  if(my_type==2 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_296.vcd");
  if(my_type==2 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_297.vcd");
  if(my_type==2 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_298.vcd");
  if(my_type==2 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_299.vcd");
  if(my_type==2 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_300.vcd");
  if(my_type==2 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_301.vcd");
  if(my_type==2 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_302.vcd");
  if(my_type==2 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_303.vcd");
  if(my_type==2 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_304.vcd");
  if(my_type==2 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_305.vcd");
  if(my_type==2 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_306.vcd");
  if(my_type==2 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_307.vcd");
  if(my_type==2 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_308.vcd");
  if(my_type==2 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_309.vcd");
  if(my_type==2 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_310.vcd");
  if(my_type==2 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_311.vcd");
  if(my_type==2 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_312.vcd");
  if(my_type==2 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_313.vcd");
  if(my_type==2 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_314.vcd");
  if(my_type==2 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_315.vcd");
  if(my_type==2 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_316.vcd");
  if(my_type==2 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_317.vcd");
  if(my_type==2 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_318.vcd");
  if(my_type==2 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_319.vcd");
  if(my_type==2 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_320.vcd");
  if(my_type==2 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_321.vcd");
  if(my_type==2 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_322.vcd");
  if(my_type==2 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_323.vcd");
  if(my_type==2 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_324.vcd");
  if(my_type==2 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_325.vcd");
  if(my_type==2 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_326.vcd");
  if(my_type==2 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_327.vcd");
  if(my_type==2 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_328.vcd");
  if(my_type==2 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_329.vcd");
  if(my_type==2 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_330.vcd");
  if(my_type==2 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_331.vcd");
  if(my_type==2 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_332.vcd");
  if(my_type==2 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_333.vcd");
  if(my_type==2 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_334.vcd");
  if(my_type==2 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_335.vcd");
  if(my_type==2 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_336.vcd");
  if(my_type==2 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_337.vcd");
  if(my_type==2 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_338.vcd");
  if(my_type==2 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_339.vcd");
  if(my_type==2 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_340.vcd");
  if(my_type==2 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_341.vcd");
  if(my_type==2 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_342.vcd");
  if(my_type==2 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_343.vcd");
  if(my_type==2 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_344.vcd");
  if(my_type==2 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_345.vcd");
  if(my_type==2 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_346.vcd");
  if(my_type==2 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_347.vcd");
  if(my_type==2 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_348.vcd");
  if(my_type==2 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_349.vcd");
  if(my_type==2 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_350.vcd");
  if(my_type==2 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_351.vcd");
  if(my_type==2 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_352.vcd");
  if(my_type==2 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_353.vcd");
  if(my_type==2 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_354.vcd");
  if(my_type==2 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_355.vcd");
  if(my_type==2 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_356.vcd");
  if(my_type==2 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_357.vcd");
  if(my_type==2 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_358.vcd");
  if(my_type==2 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_359.vcd");
  if(my_type==2 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_360.vcd");
  if(my_type==2 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_361.vcd");
  if(my_type==2 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_362.vcd");
  if(my_type==2 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_363.vcd");
  if(my_type==2 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_364.vcd");
  if(my_type==2 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_365.vcd");
  if(my_type==2 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_366.vcd");
  if(my_type==2 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_367.vcd");
  if(my_type==2 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_368.vcd");
  if(my_type==2 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_369.vcd");
  if(my_type==2 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_370.vcd");
  if(my_type==2 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_371.vcd");
  if(my_type==2 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_372.vcd");
  if(my_type==2 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_373.vcd");
  if(my_type==2 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_374.vcd");
  if(my_type==2 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_375.vcd");
  if(my_type==2 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_376.vcd");
  if(my_type==2 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_377.vcd");
  if(my_type==2 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_378.vcd");
  if(my_type==2 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_379.vcd");
  if(my_type==2 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_380.vcd");
  if(my_type==2 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_381.vcd");
  if(my_type==2 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_382.vcd");
  if(my_type==2 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_383.vcd");
  if(my_type==2 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_384.vcd");
  if(my_type==2 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_385.vcd");
  if(my_type==2 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_386.vcd");
  if(my_type==2 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_387.vcd");
  if(my_type==2 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_388.vcd");
  if(my_type==2 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_389.vcd");
  if(my_type==2 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_390.vcd");
  if(my_type==2 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_391.vcd");
  if(my_type==2 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_392.vcd");
  if(my_type==2 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_393.vcd");
  if(my_type==2 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_394.vcd");
  if(my_type==2 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_395.vcd");
  if(my_type==2 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_396.vcd");
  if(my_type==2 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_397.vcd");
  if(my_type==2 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_398.vcd");
  if(my_type==2 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_399.vcd");
  if(my_type==2 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_400.vcd");
  if(my_type==2 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_401.vcd");
  if(my_type==2 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_402.vcd");
  if(my_type==2 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_403.vcd");
  if(my_type==2 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_404.vcd");
  if(my_type==2 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_405.vcd");
  if(my_type==2 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_406.vcd");
  if(my_type==2 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_407.vcd");
  if(my_type==2 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_408.vcd");
  if(my_type==2 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_409.vcd");
  if(my_type==2 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_410.vcd");
  if(my_type==2 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_411.vcd");
  if(my_type==2 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_412.vcd");
  if(my_type==2 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_413.vcd");
  if(my_type==2 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_414.vcd");
  if(my_type==2 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_415.vcd");
  if(my_type==2 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_416.vcd");
  if(my_type==2 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_417.vcd");
  if(my_type==2 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_418.vcd");
  if(my_type==2 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_419.vcd");
  if(my_type==2 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_420.vcd");
  if(my_type==2 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_421.vcd");
  if(my_type==2 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_422.vcd");
  if(my_type==2 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_423.vcd");
  if(my_type==2 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_424.vcd");
  if(my_type==2 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_425.vcd");
  if(my_type==2 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_426.vcd");
  if(my_type==2 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_427.vcd");
  if(my_type==2 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_428.vcd");
  if(my_type==2 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_429.vcd");
  if(my_type==2 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_430.vcd");
  if(my_type==2 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_431.vcd");
  if(my_type==2 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_432.vcd");
  if(my_type==2 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_433.vcd");
  if(my_type==2 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_434.vcd");
  if(my_type==2 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_435.vcd");
  if(my_type==2 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_436.vcd");
  if(my_type==2 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_437.vcd");
  if(my_type==2 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_438.vcd");
  if(my_type==2 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_439.vcd");
  if(my_type==2 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_440.vcd");
  if(my_type==2 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_441.vcd");
  if(my_type==2 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_442.vcd");
  if(my_type==2 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_443.vcd");
  if(my_type==2 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_444.vcd");
  if(my_type==2 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_445.vcd");
  if(my_type==2 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_446.vcd");
  if(my_type==2 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_447.vcd");
  if(my_type==2 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_448.vcd");
  if(my_type==2 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_449.vcd");
  if(my_type==2 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_450.vcd");
  if(my_type==2 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_451.vcd");
  if(my_type==2 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_452.vcd");
  if(my_type==2 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_453.vcd");
  if(my_type==2 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_454.vcd");
  if(my_type==2 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_455.vcd");
  if(my_type==2 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_456.vcd");
  if(my_type==2 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_457.vcd");
  if(my_type==2 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_458.vcd");
  if(my_type==2 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_459.vcd");
  if(my_type==2 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_460.vcd");
  if(my_type==2 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_461.vcd");
  if(my_type==2 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_462.vcd");
  if(my_type==2 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_463.vcd");
  if(my_type==2 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_464.vcd");
  if(my_type==2 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_465.vcd");
  if(my_type==2 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_466.vcd");
  if(my_type==2 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_467.vcd");
  if(my_type==2 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_468.vcd");
  if(my_type==2 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_469.vcd");
  if(my_type==2 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_470.vcd");
  if(my_type==2 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_471.vcd");
  if(my_type==2 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_472.vcd");
  if(my_type==2 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_473.vcd");
  if(my_type==2 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_474.vcd");
  if(my_type==2 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_475.vcd");
  if(my_type==2 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_476.vcd");
  if(my_type==2 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_477.vcd");
  if(my_type==2 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_478.vcd");
  if(my_type==2 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_479.vcd");
  if(my_type==2 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_480.vcd");
  if(my_type==2 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_481.vcd");
  if(my_type==2 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_482.vcd");
  if(my_type==2 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_483.vcd");
  if(my_type==2 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_484.vcd");
  if(my_type==2 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_485.vcd");
  if(my_type==2 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_486.vcd");
  if(my_type==2 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_487.vcd");
  if(my_type==2 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_488.vcd");
  if(my_type==2 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_489.vcd");
  if(my_type==2 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_490.vcd");
  if(my_type==2 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_491.vcd");
  if(my_type==2 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_492.vcd");
  if(my_type==2 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_493.vcd");
  if(my_type==2 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_494.vcd");
  if(my_type==2 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_495.vcd");
  if(my_type==2 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_496.vcd");
  if(my_type==2 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_497.vcd");
  if(my_type==2 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_498.vcd");
  if(my_type==2 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_499.vcd");
  if(my_type==2 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_500.vcd");
  if(my_type==2 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_501.vcd");
  if(my_type==2 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_502.vcd");
  if(my_type==2 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_503.vcd");
  if(my_type==2 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_504.vcd");
  if(my_type==2 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_505.vcd");
  if(my_type==2 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_506.vcd");
  if(my_type==2 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_507.vcd");
  if(my_type==2 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_508.vcd");
  if(my_type==2 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_509.vcd");
  if(my_type==2 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_510.vcd");
  if(my_type==2 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_511.vcd");
  if(my_type==2 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_512.vcd");
  if(my_type==2 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_513.vcd");
  if(my_type==2 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_514.vcd");
  if(my_type==2 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_515.vcd");
  if(my_type==2 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_516.vcd");
  if(my_type==2 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_517.vcd");
  if(my_type==2 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_518.vcd");
  if(my_type==2 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_519.vcd");
  if(my_type==2 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_520.vcd");
  if(my_type==2 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_521.vcd");
  if(my_type==2 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_522.vcd");
  if(my_type==2 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_523.vcd");
  if(my_type==2 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_524.vcd");
  if(my_type==2 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_525.vcd");
  if(my_type==2 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_526.vcd");
  if(my_type==2 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_527.vcd");
  if(my_type==2 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_528.vcd");
  if(my_type==2 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_529.vcd");
  if(my_type==2 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_530.vcd");
  if(my_type==2 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_531.vcd");
  if(my_type==2 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_532.vcd");
  if(my_type==2 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_533.vcd");
  if(my_type==2 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_534.vcd");
  if(my_type==2 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_535.vcd");
  if(my_type==2 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_536.vcd");
  if(my_type==2 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_537.vcd");
  if(my_type==2 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_538.vcd");
  if(my_type==2 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_539.vcd");
  if(my_type==2 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_540.vcd");
  if(my_type==2 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_541.vcd");
  if(my_type==2 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_542.vcd");
  if(my_type==2 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_543.vcd");
  if(my_type==2 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_544.vcd");
  if(my_type==2 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_545.vcd");
  if(my_type==2 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_546.vcd");
  if(my_type==2 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_547.vcd");
  if(my_type==2 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_548.vcd");
  if(my_type==2 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_549.vcd");
  if(my_type==2 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_550.vcd");
  if(my_type==2 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_551.vcd");
  if(my_type==2 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_552.vcd");
  if(my_type==2 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_553.vcd");
  if(my_type==2 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_554.vcd");
  if(my_type==2 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_555.vcd");
  if(my_type==2 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_556.vcd");
  if(my_type==2 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_557.vcd");
  if(my_type==2 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_558.vcd");
  if(my_type==2 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_559.vcd");
  if(my_type==2 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_560.vcd");
  if(my_type==2 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_561.vcd");
  if(my_type==2 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_562.vcd");
  if(my_type==2 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_563.vcd");
  if(my_type==2 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_564.vcd");
  if(my_type==2 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_565.vcd");
  if(my_type==2 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_566.vcd");
  if(my_type==2 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_567.vcd");
  if(my_type==2 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_568.vcd");
  if(my_type==2 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_569.vcd");
  if(my_type==2 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_570.vcd");
  if(my_type==2 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_571.vcd");
  if(my_type==2 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_572.vcd");
  if(my_type==2 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_573.vcd");
  if(my_type==2 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_574.vcd");
  if(my_type==2 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_575.vcd");
  if(my_type==2 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_576.vcd");
  if(my_type==2 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_577.vcd");
  if(my_type==2 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_578.vcd");
  if(my_type==2 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_579.vcd");
  if(my_type==2 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_580.vcd");
  if(my_type==2 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_581.vcd");
  if(my_type==2 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_582.vcd");
  if(my_type==2 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_583.vcd");
  if(my_type==2 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_584.vcd");
  if(my_type==2 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_585.vcd");
  if(my_type==2 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_586.vcd");
  if(my_type==2 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_587.vcd");
  if(my_type==2 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_588.vcd");
  if(my_type==2 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_589.vcd");
  if(my_type==2 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_590.vcd");
  if(my_type==2 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_591.vcd");
  if(my_type==2 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_592.vcd");
  if(my_type==2 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_593.vcd");
  if(my_type==2 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_594.vcd");
  if(my_type==2 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_595.vcd");
  if(my_type==2 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_596.vcd");
  if(my_type==2 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_597.vcd");
  if(my_type==2 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_598.vcd");
  if(my_type==2 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_599.vcd");
  if(my_type==2 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_600.vcd");
  if(my_type==2 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_601.vcd");
  if(my_type==2 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_602.vcd");
  if(my_type==2 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_603.vcd");
  if(my_type==2 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_604.vcd");
  if(my_type==2 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_605.vcd");
  if(my_type==2 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_606.vcd");
  if(my_type==2 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_607.vcd");
  if(my_type==2 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_608.vcd");
  if(my_type==2 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_609.vcd");
  if(my_type==2 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_610.vcd");
  if(my_type==2 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_611.vcd");
  if(my_type==2 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_612.vcd");
  if(my_type==2 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_613.vcd");
  if(my_type==2 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_614.vcd");
  if(my_type==2 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_615.vcd");
  if(my_type==2 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_616.vcd");
  if(my_type==2 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_617.vcd");
  if(my_type==2 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_618.vcd");
  if(my_type==2 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_619.vcd");
  if(my_type==2 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_620.vcd");
  if(my_type==2 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_621.vcd");
  if(my_type==2 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_622.vcd");
  if(my_type==2 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_623.vcd");
  if(my_type==2 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_624.vcd");
  if(my_type==2 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_625.vcd");
  if(my_type==2 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_626.vcd");
  if(my_type==2 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_627.vcd");
  if(my_type==2 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_628.vcd");
  if(my_type==2 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_629.vcd");
  if(my_type==2 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_630.vcd");
  if(my_type==2 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_631.vcd");
  if(my_type==2 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_632.vcd");
  if(my_type==2 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_633.vcd");
  if(my_type==2 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_634.vcd");
  if(my_type==2 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_635.vcd");
  if(my_type==2 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_636.vcd");
  if(my_type==2 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_637.vcd");
  if(my_type==2 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_638.vcd");
  if(my_type==2 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_639.vcd");
  if(my_type==2 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_640.vcd");
  if(my_type==2 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_641.vcd");
  if(my_type==2 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_642.vcd");
  if(my_type==2 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_643.vcd");
  if(my_type==2 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_644.vcd");
  if(my_type==2 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_645.vcd");
  if(my_type==2 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_646.vcd");
  if(my_type==2 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_647.vcd");
  if(my_type==2 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_648.vcd");
  if(my_type==2 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_649.vcd");
  if(my_type==2 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_650.vcd");
  if(my_type==2 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_651.vcd");
  if(my_type==2 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_652.vcd");
  if(my_type==2 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_653.vcd");
  if(my_type==2 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_654.vcd");
  if(my_type==2 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_655.vcd");
  if(my_type==2 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_656.vcd");
  if(my_type==2 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_657.vcd");
  if(my_type==2 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_658.vcd");
  if(my_type==2 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_659.vcd");
  if(my_type==2 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_660.vcd");
  if(my_type==2 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_661.vcd");
  if(my_type==2 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_662.vcd");
  if(my_type==2 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_663.vcd");
  if(my_type==2 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_664.vcd");
  if(my_type==2 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_665.vcd");
  if(my_type==2 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_666.vcd");
  if(my_type==2 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_667.vcd");
  if(my_type==2 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_668.vcd");
  if(my_type==2 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_669.vcd");
  if(my_type==2 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_670.vcd");
  if(my_type==2 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_671.vcd");
  if(my_type==2 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_672.vcd");
  if(my_type==2 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_673.vcd");
  if(my_type==2 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_674.vcd");
  if(my_type==2 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_675.vcd");
  if(my_type==2 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_676.vcd");
  if(my_type==2 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_677.vcd");
  if(my_type==2 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_678.vcd");
  if(my_type==2 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_679.vcd");
  if(my_type==2 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_680.vcd");
  if(my_type==2 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_681.vcd");
  if(my_type==2 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_682.vcd");
  if(my_type==2 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_683.vcd");
  if(my_type==2 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_684.vcd");
  if(my_type==2 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_685.vcd");
  if(my_type==2 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_686.vcd");
  if(my_type==2 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_687.vcd");
  if(my_type==2 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_688.vcd");
  if(my_type==2 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_689.vcd");
  if(my_type==2 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_690.vcd");
  if(my_type==2 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_691.vcd");
  if(my_type==2 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_692.vcd");
  if(my_type==2 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_693.vcd");
  if(my_type==2 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_694.vcd");
  if(my_type==2 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_695.vcd");
  if(my_type==2 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_696.vcd");
  if(my_type==2 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_697.vcd");
  if(my_type==2 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_698.vcd");
  if(my_type==2 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_699.vcd");
  if(my_type==2 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_700.vcd");
  if(my_type==2 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_701.vcd");
  if(my_type==2 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_702.vcd");
  if(my_type==2 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_703.vcd");
  if(my_type==2 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_704.vcd");
  if(my_type==2 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_705.vcd");
  if(my_type==2 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_706.vcd");
  if(my_type==2 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_707.vcd");
  if(my_type==2 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_708.vcd");
  if(my_type==2 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_709.vcd");
  if(my_type==2 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_710.vcd");
  if(my_type==2 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_711.vcd");
  if(my_type==2 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_712.vcd");
  if(my_type==2 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_713.vcd");
  if(my_type==2 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_714.vcd");
  if(my_type==2 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_715.vcd");
  if(my_type==2 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_716.vcd");
  if(my_type==2 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_717.vcd");
  if(my_type==2 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_718.vcd");
  if(my_type==2 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_719.vcd");
  if(my_type==2 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_720.vcd");
  if(my_type==2 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_721.vcd");
  if(my_type==2 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_722.vcd");
  if(my_type==2 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_723.vcd");
  if(my_type==2 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_724.vcd");
  if(my_type==2 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_725.vcd");
  if(my_type==2 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_726.vcd");
  if(my_type==2 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_727.vcd");
  if(my_type==2 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_728.vcd");
  if(my_type==2 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_729.vcd");
  if(my_type==2 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_730.vcd");
  if(my_type==2 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_731.vcd");
  if(my_type==2 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_732.vcd");
  if(my_type==2 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_733.vcd");
  if(my_type==2 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_734.vcd");
  if(my_type==2 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_735.vcd");
  if(my_type==2 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_736.vcd");
  if(my_type==2 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_737.vcd");
  if(my_type==2 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_738.vcd");
  if(my_type==2 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_739.vcd");
  if(my_type==2 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_740.vcd");
  if(my_type==2 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_741.vcd");
  if(my_type==2 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_742.vcd");
  if(my_type==2 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_743.vcd");
  if(my_type==2 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_744.vcd");
  if(my_type==2 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_745.vcd");
  if(my_type==2 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_746.vcd");
  if(my_type==2 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_747.vcd");
  if(my_type==2 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_748.vcd");
  if(my_type==2 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_749.vcd");
  if(my_type==2 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_750.vcd");
  if(my_type==2 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_751.vcd");
  if(my_type==2 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_752.vcd");
  if(my_type==2 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_753.vcd");
  if(my_type==2 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_754.vcd");
  if(my_type==2 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_755.vcd");
  if(my_type==2 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_756.vcd");
  if(my_type==2 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_757.vcd");
  if(my_type==2 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_758.vcd");
  if(my_type==2 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_759.vcd");
  if(my_type==2 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_760.vcd");
  if(my_type==2 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_761.vcd");
  if(my_type==2 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_762.vcd");
  if(my_type==2 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_763.vcd");
  if(my_type==2 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_764.vcd");
  if(my_type==2 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_765.vcd");
  if(my_type==2 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_766.vcd");
  if(my_type==2 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_767.vcd");
  if(my_type==2 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_768.vcd");
  if(my_type==2 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_769.vcd");
  if(my_type==2 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_770.vcd");
  if(my_type==2 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_771.vcd");
  if(my_type==2 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_772.vcd");
  if(my_type==2 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_773.vcd");
  if(my_type==2 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_774.vcd");
  if(my_type==2 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_775.vcd");
  if(my_type==2 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_776.vcd");
  if(my_type==2 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_777.vcd");
  if(my_type==2 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_778.vcd");
  if(my_type==2 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_779.vcd");
  if(my_type==2 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_780.vcd");
  if(my_type==2 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_781.vcd");
  if(my_type==2 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_782.vcd");
  if(my_type==2 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_783.vcd");
  if(my_type==2 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_784.vcd");
  if(my_type==2 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_785.vcd");
  if(my_type==2 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_786.vcd");
  if(my_type==2 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_787.vcd");
  if(my_type==2 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_788.vcd");
  if(my_type==2 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_789.vcd");
  if(my_type==2 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_790.vcd");
  if(my_type==2 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_791.vcd");
  if(my_type==2 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_792.vcd");
  if(my_type==2 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_793.vcd");
  if(my_type==2 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_794.vcd");
  if(my_type==2 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_795.vcd");
  if(my_type==2 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_796.vcd");
  if(my_type==2 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_797.vcd");
  if(my_type==2 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_798.vcd");
  if(my_type==2 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_799.vcd");
  if(my_type==2 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_800.vcd");
  if(my_type==2 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_801.vcd");
  if(my_type==2 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_802.vcd");
  if(my_type==2 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_803.vcd");
  if(my_type==2 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_804.vcd");
  if(my_type==2 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_805.vcd");
  if(my_type==2 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_806.vcd");
  if(my_type==2 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_807.vcd");
  if(my_type==2 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_808.vcd");
  if(my_type==2 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_809.vcd");
  if(my_type==2 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_810.vcd");
  if(my_type==2 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_811.vcd");
  if(my_type==2 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_812.vcd");
  if(my_type==2 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_813.vcd");
  if(my_type==2 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_814.vcd");
  if(my_type==2 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_815.vcd");
  if(my_type==2 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_816.vcd");
  if(my_type==2 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_817.vcd");
  if(my_type==2 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_818.vcd");
  if(my_type==2 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_819.vcd");
  if(my_type==2 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_820.vcd");
  if(my_type==2 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_821.vcd");
  if(my_type==2 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_822.vcd");
  if(my_type==2 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_823.vcd");
  if(my_type==2 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_824.vcd");
  if(my_type==2 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_825.vcd");
  if(my_type==2 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_826.vcd");
  if(my_type==2 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_827.vcd");
  if(my_type==2 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_828.vcd");
  if(my_type==2 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_829.vcd");
  if(my_type==2 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_830.vcd");
  if(my_type==2 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_831.vcd");
  if(my_type==2 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_832.vcd");
  if(my_type==2 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_833.vcd");
  if(my_type==2 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_834.vcd");
  if(my_type==2 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_835.vcd");
  if(my_type==2 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_836.vcd");
  if(my_type==2 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_837.vcd");
  if(my_type==2 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_838.vcd");
  if(my_type==2 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_839.vcd");
  if(my_type==2 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_840.vcd");
  if(my_type==2 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_841.vcd");
  if(my_type==2 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_842.vcd");
  if(my_type==2 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_843.vcd");
  if(my_type==2 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_844.vcd");
  if(my_type==2 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_845.vcd");
  if(my_type==2 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_846.vcd");
  if(my_type==2 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_847.vcd");
  if(my_type==2 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_848.vcd");
  if(my_type==2 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_849.vcd");
  if(my_type==2 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_850.vcd");
  if(my_type==2 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_851.vcd");
  if(my_type==2 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_852.vcd");
  if(my_type==2 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_853.vcd");
  if(my_type==2 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_854.vcd");
  if(my_type==2 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_855.vcd");
  if(my_type==2 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_856.vcd");
  if(my_type==2 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_857.vcd");
  if(my_type==2 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_858.vcd");
  if(my_type==2 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_859.vcd");
  if(my_type==2 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_860.vcd");
  if(my_type==2 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_861.vcd");
  if(my_type==2 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_862.vcd");
  if(my_type==2 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_863.vcd");
  if(my_type==2 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_864.vcd");
  if(my_type==2 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_865.vcd");
  if(my_type==2 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_866.vcd");
  if(my_type==2 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_867.vcd");
  if(my_type==2 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_868.vcd");
  if(my_type==2 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_869.vcd");
  if(my_type==2 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_870.vcd");
  if(my_type==2 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_871.vcd");
  if(my_type==2 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_872.vcd");
  if(my_type==2 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_873.vcd");
  if(my_type==2 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_874.vcd");
  if(my_type==2 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_875.vcd");
  if(my_type==2 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_876.vcd");
  if(my_type==2 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_877.vcd");
  if(my_type==2 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_878.vcd");
  if(my_type==2 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_879.vcd");
  if(my_type==2 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_880.vcd");
  if(my_type==2 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_881.vcd");
  if(my_type==2 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_882.vcd");
  if(my_type==2 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_883.vcd");
  if(my_type==2 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_884.vcd");
  if(my_type==2 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_885.vcd");
  if(my_type==2 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_886.vcd");
  if(my_type==2 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_887.vcd");
  if(my_type==2 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_888.vcd");
  if(my_type==2 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_889.vcd");
  if(my_type==2 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_890.vcd");
  if(my_type==2 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_891.vcd");
  if(my_type==2 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_892.vcd");
  if(my_type==2 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_893.vcd");
  if(my_type==2 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_894.vcd");
  if(my_type==2 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_895.vcd");
  if(my_type==2 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_896.vcd");
  if(my_type==2 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_897.vcd");
  if(my_type==2 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_898.vcd");
  if(my_type==2 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_899.vcd");
  if(my_type==2 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_900.vcd");
  if(my_type==2 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_901.vcd");
  if(my_type==2 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_902.vcd");
  if(my_type==2 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_903.vcd");
  if(my_type==2 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_904.vcd");
  if(my_type==2 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_905.vcd");
  if(my_type==2 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_906.vcd");
  if(my_type==2 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_907.vcd");
  if(my_type==2 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_908.vcd");
  if(my_type==2 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_909.vcd");
  if(my_type==2 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_910.vcd");
  if(my_type==2 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_911.vcd");
  if(my_type==2 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_912.vcd");
  if(my_type==2 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_913.vcd");
  if(my_type==2 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_914.vcd");
  if(my_type==2 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_915.vcd");
  if(my_type==2 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_916.vcd");
  if(my_type==2 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_917.vcd");
  if(my_type==2 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_918.vcd");
  if(my_type==2 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_919.vcd");
  if(my_type==2 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_920.vcd");
  if(my_type==2 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_921.vcd");
  if(my_type==2 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_922.vcd");
  if(my_type==2 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_923.vcd");
  if(my_type==2 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_924.vcd");
  if(my_type==2 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_925.vcd");
  if(my_type==2 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_926.vcd");
  if(my_type==2 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_927.vcd");
  if(my_type==2 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_928.vcd");
  if(my_type==2 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_929.vcd");
  if(my_type==2 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_930.vcd");
  if(my_type==2 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_931.vcd");
  if(my_type==2 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_932.vcd");
  if(my_type==2 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_933.vcd");
  if(my_type==2 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_934.vcd");
  if(my_type==2 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_935.vcd");
  if(my_type==2 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_936.vcd");
  if(my_type==2 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_937.vcd");
  if(my_type==2 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_938.vcd");
  if(my_type==2 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_939.vcd");
  if(my_type==2 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_940.vcd");
  if(my_type==2 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_941.vcd");
  if(my_type==2 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_942.vcd");
  if(my_type==2 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_943.vcd");
  if(my_type==2 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_944.vcd");
  if(my_type==2 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_945.vcd");
  if(my_type==2 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_946.vcd");
  if(my_type==2 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_947.vcd");
  if(my_type==2 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_948.vcd");
  if(my_type==2 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_949.vcd");
  if(my_type==2 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_950.vcd");
  if(my_type==2 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_951.vcd");
  if(my_type==2 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_952.vcd");
  if(my_type==2 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_953.vcd");
  if(my_type==2 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_954.vcd");
  if(my_type==2 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_955.vcd");
  if(my_type==2 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_956.vcd");
  if(my_type==2 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_957.vcd");
  if(my_type==2 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_958.vcd");
  if(my_type==2 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_959.vcd");
  if(my_type==2 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_960.vcd");
  if(my_type==2 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_961.vcd");
  if(my_type==2 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_962.vcd");
  if(my_type==2 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_963.vcd");
  if(my_type==2 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_964.vcd");
  if(my_type==2 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_965.vcd");
  if(my_type==2 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_966.vcd");
  if(my_type==2 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_967.vcd");
  if(my_type==2 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_968.vcd");
  if(my_type==2 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_969.vcd");
  if(my_type==2 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_970.vcd");
  if(my_type==2 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_971.vcd");
  if(my_type==2 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_972.vcd");
  if(my_type==2 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_973.vcd");
  if(my_type==2 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_974.vcd");
  if(my_type==2 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_975.vcd");
  if(my_type==2 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_976.vcd");
  if(my_type==2 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_977.vcd");
  if(my_type==2 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_978.vcd");
  if(my_type==2 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_979.vcd");
  if(my_type==2 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_980.vcd");
  if(my_type==2 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_981.vcd");
  if(my_type==2 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_982.vcd");
  if(my_type==2 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_983.vcd");
  if(my_type==2 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_984.vcd");
  if(my_type==2 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_985.vcd");
  if(my_type==2 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_986.vcd");
  if(my_type==2 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_987.vcd");
  if(my_type==2 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_988.vcd");
  if(my_type==2 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_989.vcd");
  if(my_type==2 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_990.vcd");
  if(my_type==2 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_991.vcd");
  if(my_type==2 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_992.vcd");
  if(my_type==2 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_993.vcd");
  if(my_type==2 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_994.vcd");
  if(my_type==2 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_995.vcd");
  if(my_type==2 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_996.vcd");
  if(my_type==2 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_997.vcd");
  if(my_type==2 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_998.vcd");
  if(my_type==2 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_2_999.vcd");
  if(my_type==3 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_0.vcd");
  if(my_type==3 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_1.vcd");
  if(my_type==3 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_2.vcd");
  if(my_type==3 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_3.vcd");
  if(my_type==3 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_4.vcd");
  if(my_type==3 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_5.vcd");
  if(my_type==3 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_6.vcd");
  if(my_type==3 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_7.vcd");
  if(my_type==3 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_8.vcd");
  if(my_type==3 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_9.vcd");
  if(my_type==3 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_10.vcd");
  if(my_type==3 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_11.vcd");
  if(my_type==3 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_12.vcd");
  if(my_type==3 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_13.vcd");
  if(my_type==3 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_14.vcd");
  if(my_type==3 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_15.vcd");
  if(my_type==3 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_16.vcd");
  if(my_type==3 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_17.vcd");
  if(my_type==3 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_18.vcd");
  if(my_type==3 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_19.vcd");
  if(my_type==3 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_20.vcd");
  if(my_type==3 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_21.vcd");
  if(my_type==3 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_22.vcd");
  if(my_type==3 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_23.vcd");
  if(my_type==3 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_24.vcd");
  if(my_type==3 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_25.vcd");
  if(my_type==3 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_26.vcd");
  if(my_type==3 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_27.vcd");
  if(my_type==3 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_28.vcd");
  if(my_type==3 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_29.vcd");
  if(my_type==3 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_30.vcd");
  if(my_type==3 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_31.vcd");
  if(my_type==3 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_32.vcd");
  if(my_type==3 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_33.vcd");
  if(my_type==3 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_34.vcd");
  if(my_type==3 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_35.vcd");
  if(my_type==3 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_36.vcd");
  if(my_type==3 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_37.vcd");
  if(my_type==3 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_38.vcd");
  if(my_type==3 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_39.vcd");
  if(my_type==3 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_40.vcd");
  if(my_type==3 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_41.vcd");
  if(my_type==3 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_42.vcd");
  if(my_type==3 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_43.vcd");
  if(my_type==3 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_44.vcd");
  if(my_type==3 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_45.vcd");
  if(my_type==3 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_46.vcd");
  if(my_type==3 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_47.vcd");
  if(my_type==3 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_48.vcd");
  if(my_type==3 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_49.vcd");
  if(my_type==3 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_50.vcd");
  if(my_type==3 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_51.vcd");
  if(my_type==3 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_52.vcd");
  if(my_type==3 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_53.vcd");
  if(my_type==3 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_54.vcd");
  if(my_type==3 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_55.vcd");
  if(my_type==3 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_56.vcd");
  if(my_type==3 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_57.vcd");
  if(my_type==3 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_58.vcd");
  if(my_type==3 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_59.vcd");
  if(my_type==3 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_60.vcd");
  if(my_type==3 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_61.vcd");
  if(my_type==3 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_62.vcd");
  if(my_type==3 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_63.vcd");
  if(my_type==3 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_64.vcd");
  if(my_type==3 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_65.vcd");
  if(my_type==3 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_66.vcd");
  if(my_type==3 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_67.vcd");
  if(my_type==3 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_68.vcd");
  if(my_type==3 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_69.vcd");
  if(my_type==3 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_70.vcd");
  if(my_type==3 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_71.vcd");
  if(my_type==3 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_72.vcd");
  if(my_type==3 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_73.vcd");
  if(my_type==3 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_74.vcd");
  if(my_type==3 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_75.vcd");
  if(my_type==3 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_76.vcd");
  if(my_type==3 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_77.vcd");
  if(my_type==3 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_78.vcd");
  if(my_type==3 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_79.vcd");
  if(my_type==3 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_80.vcd");
  if(my_type==3 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_81.vcd");
  if(my_type==3 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_82.vcd");
  if(my_type==3 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_83.vcd");
  if(my_type==3 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_84.vcd");
  if(my_type==3 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_85.vcd");
  if(my_type==3 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_86.vcd");
  if(my_type==3 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_87.vcd");
  if(my_type==3 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_88.vcd");
  if(my_type==3 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_89.vcd");
  if(my_type==3 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_90.vcd");
  if(my_type==3 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_91.vcd");
  if(my_type==3 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_92.vcd");
  if(my_type==3 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_93.vcd");
  if(my_type==3 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_94.vcd");
  if(my_type==3 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_95.vcd");
  if(my_type==3 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_96.vcd");
  if(my_type==3 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_97.vcd");
  if(my_type==3 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_98.vcd");
  if(my_type==3 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_99.vcd");
  if(my_type==3 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_100.vcd");
  if(my_type==3 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_101.vcd");
  if(my_type==3 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_102.vcd");
  if(my_type==3 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_103.vcd");
  if(my_type==3 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_104.vcd");
  if(my_type==3 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_105.vcd");
  if(my_type==3 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_106.vcd");
  if(my_type==3 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_107.vcd");
  if(my_type==3 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_108.vcd");
  if(my_type==3 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_109.vcd");
  if(my_type==3 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_110.vcd");
  if(my_type==3 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_111.vcd");
  if(my_type==3 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_112.vcd");
  if(my_type==3 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_113.vcd");
  if(my_type==3 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_114.vcd");
  if(my_type==3 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_115.vcd");
  if(my_type==3 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_116.vcd");
  if(my_type==3 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_117.vcd");
  if(my_type==3 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_118.vcd");
  if(my_type==3 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_119.vcd");
  if(my_type==3 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_120.vcd");
  if(my_type==3 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_121.vcd");
  if(my_type==3 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_122.vcd");
  if(my_type==3 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_123.vcd");
  if(my_type==3 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_124.vcd");
  if(my_type==3 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_125.vcd");
  if(my_type==3 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_126.vcd");
  if(my_type==3 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_127.vcd");
  if(my_type==3 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_128.vcd");
  if(my_type==3 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_129.vcd");
  if(my_type==3 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_130.vcd");
  if(my_type==3 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_131.vcd");
  if(my_type==3 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_132.vcd");
  if(my_type==3 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_133.vcd");
  if(my_type==3 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_134.vcd");
  if(my_type==3 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_135.vcd");
  if(my_type==3 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_136.vcd");
  if(my_type==3 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_137.vcd");
  if(my_type==3 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_138.vcd");
  if(my_type==3 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_139.vcd");
  if(my_type==3 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_140.vcd");
  if(my_type==3 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_141.vcd");
  if(my_type==3 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_142.vcd");
  if(my_type==3 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_143.vcd");
  if(my_type==3 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_144.vcd");
  if(my_type==3 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_145.vcd");
  if(my_type==3 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_146.vcd");
  if(my_type==3 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_147.vcd");
  if(my_type==3 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_148.vcd");
  if(my_type==3 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_149.vcd");
  if(my_type==3 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_150.vcd");
  if(my_type==3 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_151.vcd");
  if(my_type==3 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_152.vcd");
  if(my_type==3 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_153.vcd");
  if(my_type==3 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_154.vcd");
  if(my_type==3 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_155.vcd");
  if(my_type==3 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_156.vcd");
  if(my_type==3 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_157.vcd");
  if(my_type==3 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_158.vcd");
  if(my_type==3 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_159.vcd");
  if(my_type==3 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_160.vcd");
  if(my_type==3 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_161.vcd");
  if(my_type==3 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_162.vcd");
  if(my_type==3 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_163.vcd");
  if(my_type==3 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_164.vcd");
  if(my_type==3 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_165.vcd");
  if(my_type==3 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_166.vcd");
  if(my_type==3 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_167.vcd");
  if(my_type==3 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_168.vcd");
  if(my_type==3 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_169.vcd");
  if(my_type==3 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_170.vcd");
  if(my_type==3 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_171.vcd");
  if(my_type==3 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_172.vcd");
  if(my_type==3 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_173.vcd");
  if(my_type==3 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_174.vcd");
  if(my_type==3 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_175.vcd");
  if(my_type==3 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_176.vcd");
  if(my_type==3 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_177.vcd");
  if(my_type==3 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_178.vcd");
  if(my_type==3 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_179.vcd");
  if(my_type==3 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_180.vcd");
  if(my_type==3 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_181.vcd");
  if(my_type==3 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_182.vcd");
  if(my_type==3 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_183.vcd");
  if(my_type==3 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_184.vcd");
  if(my_type==3 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_185.vcd");
  if(my_type==3 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_186.vcd");
  if(my_type==3 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_187.vcd");
  if(my_type==3 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_188.vcd");
  if(my_type==3 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_189.vcd");
  if(my_type==3 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_190.vcd");
  if(my_type==3 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_191.vcd");
  if(my_type==3 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_192.vcd");
  if(my_type==3 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_193.vcd");
  if(my_type==3 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_194.vcd");
  if(my_type==3 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_195.vcd");
  if(my_type==3 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_196.vcd");
  if(my_type==3 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_197.vcd");
  if(my_type==3 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_198.vcd");
  if(my_type==3 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_199.vcd");
  if(my_type==3 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_200.vcd");
  if(my_type==3 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_201.vcd");
  if(my_type==3 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_202.vcd");
  if(my_type==3 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_203.vcd");
  if(my_type==3 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_204.vcd");
  if(my_type==3 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_205.vcd");
  if(my_type==3 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_206.vcd");
  if(my_type==3 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_207.vcd");
  if(my_type==3 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_208.vcd");
  if(my_type==3 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_209.vcd");
  if(my_type==3 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_210.vcd");
  if(my_type==3 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_211.vcd");
  if(my_type==3 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_212.vcd");
  if(my_type==3 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_213.vcd");
  if(my_type==3 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_214.vcd");
  if(my_type==3 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_215.vcd");
  if(my_type==3 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_216.vcd");
  if(my_type==3 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_217.vcd");
  if(my_type==3 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_218.vcd");
  if(my_type==3 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_219.vcd");
  if(my_type==3 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_220.vcd");
  if(my_type==3 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_221.vcd");
  if(my_type==3 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_222.vcd");
  if(my_type==3 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_223.vcd");
  if(my_type==3 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_224.vcd");
  if(my_type==3 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_225.vcd");
  if(my_type==3 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_226.vcd");
  if(my_type==3 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_227.vcd");
  if(my_type==3 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_228.vcd");
  if(my_type==3 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_229.vcd");
  if(my_type==3 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_230.vcd");
  if(my_type==3 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_231.vcd");
  if(my_type==3 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_232.vcd");
  if(my_type==3 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_233.vcd");
  if(my_type==3 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_234.vcd");
  if(my_type==3 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_235.vcd");
  if(my_type==3 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_236.vcd");
  if(my_type==3 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_237.vcd");
  if(my_type==3 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_238.vcd");
  if(my_type==3 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_239.vcd");
  if(my_type==3 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_240.vcd");
  if(my_type==3 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_241.vcd");
  if(my_type==3 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_242.vcd");
  if(my_type==3 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_243.vcd");
  if(my_type==3 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_244.vcd");
  if(my_type==3 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_245.vcd");
  if(my_type==3 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_246.vcd");
  if(my_type==3 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_247.vcd");
  if(my_type==3 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_248.vcd");
  if(my_type==3 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_249.vcd");
  if(my_type==3 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_250.vcd");
  if(my_type==3 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_251.vcd");
  if(my_type==3 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_252.vcd");
  if(my_type==3 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_253.vcd");
  if(my_type==3 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_254.vcd");
  if(my_type==3 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_255.vcd");
  if(my_type==3 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_256.vcd");
  if(my_type==3 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_257.vcd");
  if(my_type==3 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_258.vcd");
  if(my_type==3 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_259.vcd");
  if(my_type==3 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_260.vcd");
  if(my_type==3 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_261.vcd");
  if(my_type==3 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_262.vcd");
  if(my_type==3 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_263.vcd");
  if(my_type==3 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_264.vcd");
  if(my_type==3 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_265.vcd");
  if(my_type==3 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_266.vcd");
  if(my_type==3 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_267.vcd");
  if(my_type==3 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_268.vcd");
  if(my_type==3 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_269.vcd");
  if(my_type==3 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_270.vcd");
  if(my_type==3 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_271.vcd");
  if(my_type==3 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_272.vcd");
  if(my_type==3 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_273.vcd");
  if(my_type==3 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_274.vcd");
  if(my_type==3 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_275.vcd");
  if(my_type==3 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_276.vcd");
  if(my_type==3 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_277.vcd");
  if(my_type==3 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_278.vcd");
  if(my_type==3 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_279.vcd");
  if(my_type==3 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_280.vcd");
  if(my_type==3 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_281.vcd");
  if(my_type==3 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_282.vcd");
  if(my_type==3 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_283.vcd");
  if(my_type==3 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_284.vcd");
  if(my_type==3 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_285.vcd");
  if(my_type==3 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_286.vcd");
  if(my_type==3 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_287.vcd");
  if(my_type==3 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_288.vcd");
  if(my_type==3 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_289.vcd");
  if(my_type==3 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_290.vcd");
  if(my_type==3 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_291.vcd");
  if(my_type==3 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_292.vcd");
  if(my_type==3 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_293.vcd");
  if(my_type==3 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_294.vcd");
  if(my_type==3 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_295.vcd");
  if(my_type==3 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_296.vcd");
  if(my_type==3 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_297.vcd");
  if(my_type==3 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_298.vcd");
  if(my_type==3 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_299.vcd");
  if(my_type==3 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_300.vcd");
  if(my_type==3 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_301.vcd");
  if(my_type==3 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_302.vcd");
  if(my_type==3 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_303.vcd");
  if(my_type==3 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_304.vcd");
  if(my_type==3 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_305.vcd");
  if(my_type==3 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_306.vcd");
  if(my_type==3 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_307.vcd");
  if(my_type==3 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_308.vcd");
  if(my_type==3 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_309.vcd");
  if(my_type==3 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_310.vcd");
  if(my_type==3 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_311.vcd");
  if(my_type==3 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_312.vcd");
  if(my_type==3 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_313.vcd");
  if(my_type==3 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_314.vcd");
  if(my_type==3 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_315.vcd");
  if(my_type==3 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_316.vcd");
  if(my_type==3 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_317.vcd");
  if(my_type==3 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_318.vcd");
  if(my_type==3 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_319.vcd");
  if(my_type==3 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_320.vcd");
  if(my_type==3 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_321.vcd");
  if(my_type==3 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_322.vcd");
  if(my_type==3 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_323.vcd");
  if(my_type==3 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_324.vcd");
  if(my_type==3 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_325.vcd");
  if(my_type==3 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_326.vcd");
  if(my_type==3 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_327.vcd");
  if(my_type==3 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_328.vcd");
  if(my_type==3 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_329.vcd");
  if(my_type==3 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_330.vcd");
  if(my_type==3 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_331.vcd");
  if(my_type==3 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_332.vcd");
  if(my_type==3 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_333.vcd");
  if(my_type==3 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_334.vcd");
  if(my_type==3 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_335.vcd");
  if(my_type==3 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_336.vcd");
  if(my_type==3 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_337.vcd");
  if(my_type==3 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_338.vcd");
  if(my_type==3 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_339.vcd");
  if(my_type==3 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_340.vcd");
  if(my_type==3 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_341.vcd");
  if(my_type==3 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_342.vcd");
  if(my_type==3 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_343.vcd");
  if(my_type==3 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_344.vcd");
  if(my_type==3 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_345.vcd");
  if(my_type==3 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_346.vcd");
  if(my_type==3 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_347.vcd");
  if(my_type==3 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_348.vcd");
  if(my_type==3 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_349.vcd");
  if(my_type==3 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_350.vcd");
  if(my_type==3 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_351.vcd");
  if(my_type==3 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_352.vcd");
  if(my_type==3 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_353.vcd");
  if(my_type==3 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_354.vcd");
  if(my_type==3 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_355.vcd");
  if(my_type==3 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_356.vcd");
  if(my_type==3 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_357.vcd");
  if(my_type==3 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_358.vcd");
  if(my_type==3 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_359.vcd");
  if(my_type==3 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_360.vcd");
  if(my_type==3 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_361.vcd");
  if(my_type==3 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_362.vcd");
  if(my_type==3 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_363.vcd");
  if(my_type==3 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_364.vcd");
  if(my_type==3 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_365.vcd");
  if(my_type==3 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_366.vcd");
  if(my_type==3 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_367.vcd");
  if(my_type==3 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_368.vcd");
  if(my_type==3 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_369.vcd");
  if(my_type==3 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_370.vcd");
  if(my_type==3 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_371.vcd");
  if(my_type==3 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_372.vcd");
  if(my_type==3 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_373.vcd");
  if(my_type==3 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_374.vcd");
  if(my_type==3 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_375.vcd");
  if(my_type==3 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_376.vcd");
  if(my_type==3 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_377.vcd");
  if(my_type==3 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_378.vcd");
  if(my_type==3 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_379.vcd");
  if(my_type==3 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_380.vcd");
  if(my_type==3 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_381.vcd");
  if(my_type==3 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_382.vcd");
  if(my_type==3 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_383.vcd");
  if(my_type==3 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_384.vcd");
  if(my_type==3 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_385.vcd");
  if(my_type==3 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_386.vcd");
  if(my_type==3 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_387.vcd");
  if(my_type==3 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_388.vcd");
  if(my_type==3 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_389.vcd");
  if(my_type==3 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_390.vcd");
  if(my_type==3 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_391.vcd");
  if(my_type==3 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_392.vcd");
  if(my_type==3 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_393.vcd");
  if(my_type==3 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_394.vcd");
  if(my_type==3 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_395.vcd");
  if(my_type==3 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_396.vcd");
  if(my_type==3 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_397.vcd");
  if(my_type==3 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_398.vcd");
  if(my_type==3 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_399.vcd");
  if(my_type==3 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_400.vcd");
  if(my_type==3 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_401.vcd");
  if(my_type==3 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_402.vcd");
  if(my_type==3 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_403.vcd");
  if(my_type==3 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_404.vcd");
  if(my_type==3 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_405.vcd");
  if(my_type==3 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_406.vcd");
  if(my_type==3 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_407.vcd");
  if(my_type==3 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_408.vcd");
  if(my_type==3 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_409.vcd");
  if(my_type==3 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_410.vcd");
  if(my_type==3 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_411.vcd");
  if(my_type==3 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_412.vcd");
  if(my_type==3 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_413.vcd");
  if(my_type==3 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_414.vcd");
  if(my_type==3 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_415.vcd");
  if(my_type==3 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_416.vcd");
  if(my_type==3 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_417.vcd");
  if(my_type==3 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_418.vcd");
  if(my_type==3 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_419.vcd");
  if(my_type==3 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_420.vcd");
  if(my_type==3 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_421.vcd");
  if(my_type==3 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_422.vcd");
  if(my_type==3 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_423.vcd");
  if(my_type==3 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_424.vcd");
  if(my_type==3 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_425.vcd");
  if(my_type==3 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_426.vcd");
  if(my_type==3 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_427.vcd");
  if(my_type==3 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_428.vcd");
  if(my_type==3 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_429.vcd");
  if(my_type==3 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_430.vcd");
  if(my_type==3 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_431.vcd");
  if(my_type==3 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_432.vcd");
  if(my_type==3 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_433.vcd");
  if(my_type==3 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_434.vcd");
  if(my_type==3 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_435.vcd");
  if(my_type==3 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_436.vcd");
  if(my_type==3 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_437.vcd");
  if(my_type==3 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_438.vcd");
  if(my_type==3 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_439.vcd");
  if(my_type==3 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_440.vcd");
  if(my_type==3 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_441.vcd");
  if(my_type==3 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_442.vcd");
  if(my_type==3 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_443.vcd");
  if(my_type==3 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_444.vcd");
  if(my_type==3 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_445.vcd");
  if(my_type==3 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_446.vcd");
  if(my_type==3 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_447.vcd");
  if(my_type==3 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_448.vcd");
  if(my_type==3 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_449.vcd");
  if(my_type==3 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_450.vcd");
  if(my_type==3 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_451.vcd");
  if(my_type==3 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_452.vcd");
  if(my_type==3 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_453.vcd");
  if(my_type==3 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_454.vcd");
  if(my_type==3 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_455.vcd");
  if(my_type==3 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_456.vcd");
  if(my_type==3 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_457.vcd");
  if(my_type==3 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_458.vcd");
  if(my_type==3 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_459.vcd");
  if(my_type==3 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_460.vcd");
  if(my_type==3 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_461.vcd");
  if(my_type==3 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_462.vcd");
  if(my_type==3 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_463.vcd");
  if(my_type==3 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_464.vcd");
  if(my_type==3 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_465.vcd");
  if(my_type==3 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_466.vcd");
  if(my_type==3 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_467.vcd");
  if(my_type==3 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_468.vcd");
  if(my_type==3 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_469.vcd");
  if(my_type==3 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_470.vcd");
  if(my_type==3 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_471.vcd");
  if(my_type==3 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_472.vcd");
  if(my_type==3 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_473.vcd");
  if(my_type==3 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_474.vcd");
  if(my_type==3 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_475.vcd");
  if(my_type==3 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_476.vcd");
  if(my_type==3 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_477.vcd");
  if(my_type==3 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_478.vcd");
  if(my_type==3 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_479.vcd");
  if(my_type==3 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_480.vcd");
  if(my_type==3 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_481.vcd");
  if(my_type==3 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_482.vcd");
  if(my_type==3 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_483.vcd");
  if(my_type==3 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_484.vcd");
  if(my_type==3 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_485.vcd");
  if(my_type==3 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_486.vcd");
  if(my_type==3 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_487.vcd");
  if(my_type==3 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_488.vcd");
  if(my_type==3 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_489.vcd");
  if(my_type==3 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_490.vcd");
  if(my_type==3 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_491.vcd");
  if(my_type==3 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_492.vcd");
  if(my_type==3 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_493.vcd");
  if(my_type==3 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_494.vcd");
  if(my_type==3 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_495.vcd");
  if(my_type==3 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_496.vcd");
  if(my_type==3 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_497.vcd");
  if(my_type==3 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_498.vcd");
  if(my_type==3 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_499.vcd");
  if(my_type==3 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_500.vcd");
  if(my_type==3 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_501.vcd");
  if(my_type==3 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_502.vcd");
  if(my_type==3 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_503.vcd");
  if(my_type==3 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_504.vcd");
  if(my_type==3 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_505.vcd");
  if(my_type==3 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_506.vcd");
  if(my_type==3 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_507.vcd");
  if(my_type==3 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_508.vcd");
  if(my_type==3 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_509.vcd");
  if(my_type==3 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_510.vcd");
  if(my_type==3 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_511.vcd");
  if(my_type==3 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_512.vcd");
  if(my_type==3 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_513.vcd");
  if(my_type==3 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_514.vcd");
  if(my_type==3 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_515.vcd");
  if(my_type==3 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_516.vcd");
  if(my_type==3 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_517.vcd");
  if(my_type==3 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_518.vcd");
  if(my_type==3 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_519.vcd");
  if(my_type==3 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_520.vcd");
  if(my_type==3 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_521.vcd");
  if(my_type==3 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_522.vcd");
  if(my_type==3 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_523.vcd");
  if(my_type==3 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_524.vcd");
  if(my_type==3 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_525.vcd");
  if(my_type==3 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_526.vcd");
  if(my_type==3 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_527.vcd");
  if(my_type==3 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_528.vcd");
  if(my_type==3 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_529.vcd");
  if(my_type==3 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_530.vcd");
  if(my_type==3 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_531.vcd");
  if(my_type==3 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_532.vcd");
  if(my_type==3 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_533.vcd");
  if(my_type==3 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_534.vcd");
  if(my_type==3 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_535.vcd");
  if(my_type==3 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_536.vcd");
  if(my_type==3 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_537.vcd");
  if(my_type==3 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_538.vcd");
  if(my_type==3 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_539.vcd");
  if(my_type==3 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_540.vcd");
  if(my_type==3 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_541.vcd");
  if(my_type==3 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_542.vcd");
  if(my_type==3 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_543.vcd");
  if(my_type==3 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_544.vcd");
  if(my_type==3 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_545.vcd");
  if(my_type==3 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_546.vcd");
  if(my_type==3 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_547.vcd");
  if(my_type==3 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_548.vcd");
  if(my_type==3 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_549.vcd");
  if(my_type==3 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_550.vcd");
  if(my_type==3 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_551.vcd");
  if(my_type==3 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_552.vcd");
  if(my_type==3 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_553.vcd");
  if(my_type==3 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_554.vcd");
  if(my_type==3 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_555.vcd");
  if(my_type==3 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_556.vcd");
  if(my_type==3 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_557.vcd");
  if(my_type==3 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_558.vcd");
  if(my_type==3 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_559.vcd");
  if(my_type==3 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_560.vcd");
  if(my_type==3 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_561.vcd");
  if(my_type==3 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_562.vcd");
  if(my_type==3 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_563.vcd");
  if(my_type==3 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_564.vcd");
  if(my_type==3 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_565.vcd");
  if(my_type==3 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_566.vcd");
  if(my_type==3 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_567.vcd");
  if(my_type==3 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_568.vcd");
  if(my_type==3 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_569.vcd");
  if(my_type==3 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_570.vcd");
  if(my_type==3 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_571.vcd");
  if(my_type==3 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_572.vcd");
  if(my_type==3 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_573.vcd");
  if(my_type==3 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_574.vcd");
  if(my_type==3 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_575.vcd");
  if(my_type==3 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_576.vcd");
  if(my_type==3 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_577.vcd");
  if(my_type==3 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_578.vcd");
  if(my_type==3 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_579.vcd");
  if(my_type==3 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_580.vcd");
  if(my_type==3 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_581.vcd");
  if(my_type==3 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_582.vcd");
  if(my_type==3 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_583.vcd");
  if(my_type==3 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_584.vcd");
  if(my_type==3 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_585.vcd");
  if(my_type==3 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_586.vcd");
  if(my_type==3 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_587.vcd");
  if(my_type==3 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_588.vcd");
  if(my_type==3 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_589.vcd");
  if(my_type==3 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_590.vcd");
  if(my_type==3 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_591.vcd");
  if(my_type==3 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_592.vcd");
  if(my_type==3 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_593.vcd");
  if(my_type==3 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_594.vcd");
  if(my_type==3 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_595.vcd");
  if(my_type==3 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_596.vcd");
  if(my_type==3 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_597.vcd");
  if(my_type==3 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_598.vcd");
  if(my_type==3 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_599.vcd");
  if(my_type==3 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_600.vcd");
  if(my_type==3 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_601.vcd");
  if(my_type==3 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_602.vcd");
  if(my_type==3 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_603.vcd");
  if(my_type==3 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_604.vcd");
  if(my_type==3 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_605.vcd");
  if(my_type==3 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_606.vcd");
  if(my_type==3 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_607.vcd");
  if(my_type==3 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_608.vcd");
  if(my_type==3 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_609.vcd");
  if(my_type==3 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_610.vcd");
  if(my_type==3 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_611.vcd");
  if(my_type==3 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_612.vcd");
  if(my_type==3 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_613.vcd");
  if(my_type==3 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_614.vcd");
  if(my_type==3 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_615.vcd");
  if(my_type==3 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_616.vcd");
  if(my_type==3 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_617.vcd");
  if(my_type==3 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_618.vcd");
  if(my_type==3 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_619.vcd");
  if(my_type==3 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_620.vcd");
  if(my_type==3 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_621.vcd");
  if(my_type==3 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_622.vcd");
  if(my_type==3 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_623.vcd");
  if(my_type==3 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_624.vcd");
  if(my_type==3 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_625.vcd");
  if(my_type==3 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_626.vcd");
  if(my_type==3 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_627.vcd");
  if(my_type==3 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_628.vcd");
  if(my_type==3 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_629.vcd");
  if(my_type==3 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_630.vcd");
  if(my_type==3 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_631.vcd");
  if(my_type==3 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_632.vcd");
  if(my_type==3 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_633.vcd");
  if(my_type==3 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_634.vcd");
  if(my_type==3 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_635.vcd");
  if(my_type==3 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_636.vcd");
  if(my_type==3 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_637.vcd");
  if(my_type==3 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_638.vcd");
  if(my_type==3 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_639.vcd");
  if(my_type==3 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_640.vcd");
  if(my_type==3 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_641.vcd");
  if(my_type==3 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_642.vcd");
  if(my_type==3 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_643.vcd");
  if(my_type==3 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_644.vcd");
  if(my_type==3 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_645.vcd");
  if(my_type==3 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_646.vcd");
  if(my_type==3 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_647.vcd");
  if(my_type==3 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_648.vcd");
  if(my_type==3 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_649.vcd");
  if(my_type==3 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_650.vcd");
  if(my_type==3 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_651.vcd");
  if(my_type==3 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_652.vcd");
  if(my_type==3 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_653.vcd");
  if(my_type==3 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_654.vcd");
  if(my_type==3 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_655.vcd");
  if(my_type==3 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_656.vcd");
  if(my_type==3 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_657.vcd");
  if(my_type==3 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_658.vcd");
  if(my_type==3 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_659.vcd");
  if(my_type==3 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_660.vcd");
  if(my_type==3 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_661.vcd");
  if(my_type==3 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_662.vcd");
  if(my_type==3 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_663.vcd");
  if(my_type==3 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_664.vcd");
  if(my_type==3 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_665.vcd");
  if(my_type==3 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_666.vcd");
  if(my_type==3 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_667.vcd");
  if(my_type==3 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_668.vcd");
  if(my_type==3 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_669.vcd");
  if(my_type==3 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_670.vcd");
  if(my_type==3 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_671.vcd");
  if(my_type==3 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_672.vcd");
  if(my_type==3 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_673.vcd");
  if(my_type==3 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_674.vcd");
  if(my_type==3 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_675.vcd");
  if(my_type==3 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_676.vcd");
  if(my_type==3 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_677.vcd");
  if(my_type==3 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_678.vcd");
  if(my_type==3 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_679.vcd");
  if(my_type==3 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_680.vcd");
  if(my_type==3 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_681.vcd");
  if(my_type==3 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_682.vcd");
  if(my_type==3 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_683.vcd");
  if(my_type==3 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_684.vcd");
  if(my_type==3 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_685.vcd");
  if(my_type==3 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_686.vcd");
  if(my_type==3 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_687.vcd");
  if(my_type==3 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_688.vcd");
  if(my_type==3 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_689.vcd");
  if(my_type==3 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_690.vcd");
  if(my_type==3 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_691.vcd");
  if(my_type==3 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_692.vcd");
  if(my_type==3 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_693.vcd");
  if(my_type==3 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_694.vcd");
  if(my_type==3 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_695.vcd");
  if(my_type==3 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_696.vcd");
  if(my_type==3 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_697.vcd");
  if(my_type==3 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_698.vcd");
  if(my_type==3 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_699.vcd");
  if(my_type==3 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_700.vcd");
  if(my_type==3 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_701.vcd");
  if(my_type==3 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_702.vcd");
  if(my_type==3 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_703.vcd");
  if(my_type==3 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_704.vcd");
  if(my_type==3 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_705.vcd");
  if(my_type==3 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_706.vcd");
  if(my_type==3 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_707.vcd");
  if(my_type==3 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_708.vcd");
  if(my_type==3 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_709.vcd");
  if(my_type==3 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_710.vcd");
  if(my_type==3 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_711.vcd");
  if(my_type==3 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_712.vcd");
  if(my_type==3 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_713.vcd");
  if(my_type==3 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_714.vcd");
  if(my_type==3 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_715.vcd");
  if(my_type==3 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_716.vcd");
  if(my_type==3 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_717.vcd");
  if(my_type==3 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_718.vcd");
  if(my_type==3 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_719.vcd");
  if(my_type==3 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_720.vcd");
  if(my_type==3 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_721.vcd");
  if(my_type==3 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_722.vcd");
  if(my_type==3 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_723.vcd");
  if(my_type==3 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_724.vcd");
  if(my_type==3 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_725.vcd");
  if(my_type==3 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_726.vcd");
  if(my_type==3 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_727.vcd");
  if(my_type==3 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_728.vcd");
  if(my_type==3 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_729.vcd");
  if(my_type==3 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_730.vcd");
  if(my_type==3 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_731.vcd");
  if(my_type==3 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_732.vcd");
  if(my_type==3 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_733.vcd");
  if(my_type==3 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_734.vcd");
  if(my_type==3 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_735.vcd");
  if(my_type==3 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_736.vcd");
  if(my_type==3 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_737.vcd");
  if(my_type==3 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_738.vcd");
  if(my_type==3 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_739.vcd");
  if(my_type==3 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_740.vcd");
  if(my_type==3 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_741.vcd");
  if(my_type==3 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_742.vcd");
  if(my_type==3 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_743.vcd");
  if(my_type==3 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_744.vcd");
  if(my_type==3 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_745.vcd");
  if(my_type==3 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_746.vcd");
  if(my_type==3 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_747.vcd");
  if(my_type==3 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_748.vcd");
  if(my_type==3 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_749.vcd");
  if(my_type==3 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_750.vcd");
  if(my_type==3 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_751.vcd");
  if(my_type==3 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_752.vcd");
  if(my_type==3 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_753.vcd");
  if(my_type==3 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_754.vcd");
  if(my_type==3 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_755.vcd");
  if(my_type==3 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_756.vcd");
  if(my_type==3 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_757.vcd");
  if(my_type==3 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_758.vcd");
  if(my_type==3 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_759.vcd");
  if(my_type==3 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_760.vcd");
  if(my_type==3 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_761.vcd");
  if(my_type==3 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_762.vcd");
  if(my_type==3 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_763.vcd");
  if(my_type==3 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_764.vcd");
  if(my_type==3 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_765.vcd");
  if(my_type==3 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_766.vcd");
  if(my_type==3 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_767.vcd");
  if(my_type==3 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_768.vcd");
  if(my_type==3 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_769.vcd");
  if(my_type==3 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_770.vcd");
  if(my_type==3 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_771.vcd");
  if(my_type==3 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_772.vcd");
  if(my_type==3 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_773.vcd");
  if(my_type==3 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_774.vcd");
  if(my_type==3 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_775.vcd");
  if(my_type==3 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_776.vcd");
  if(my_type==3 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_777.vcd");
  if(my_type==3 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_778.vcd");
  if(my_type==3 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_779.vcd");
  if(my_type==3 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_780.vcd");
  if(my_type==3 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_781.vcd");
  if(my_type==3 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_782.vcd");
  if(my_type==3 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_783.vcd");
  if(my_type==3 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_784.vcd");
  if(my_type==3 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_785.vcd");
  if(my_type==3 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_786.vcd");
  if(my_type==3 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_787.vcd");
  if(my_type==3 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_788.vcd");
  if(my_type==3 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_789.vcd");
  if(my_type==3 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_790.vcd");
  if(my_type==3 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_791.vcd");
  if(my_type==3 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_792.vcd");
  if(my_type==3 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_793.vcd");
  if(my_type==3 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_794.vcd");
  if(my_type==3 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_795.vcd");
  if(my_type==3 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_796.vcd");
  if(my_type==3 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_797.vcd");
  if(my_type==3 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_798.vcd");
  if(my_type==3 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_799.vcd");
  if(my_type==3 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_800.vcd");
  if(my_type==3 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_801.vcd");
  if(my_type==3 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_802.vcd");
  if(my_type==3 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_803.vcd");
  if(my_type==3 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_804.vcd");
  if(my_type==3 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_805.vcd");
  if(my_type==3 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_806.vcd");
  if(my_type==3 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_807.vcd");
  if(my_type==3 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_808.vcd");
  if(my_type==3 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_809.vcd");
  if(my_type==3 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_810.vcd");
  if(my_type==3 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_811.vcd");
  if(my_type==3 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_812.vcd");
  if(my_type==3 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_813.vcd");
  if(my_type==3 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_814.vcd");
  if(my_type==3 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_815.vcd");
  if(my_type==3 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_816.vcd");
  if(my_type==3 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_817.vcd");
  if(my_type==3 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_818.vcd");
  if(my_type==3 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_819.vcd");
  if(my_type==3 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_820.vcd");
  if(my_type==3 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_821.vcd");
  if(my_type==3 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_822.vcd");
  if(my_type==3 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_823.vcd");
  if(my_type==3 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_824.vcd");
  if(my_type==3 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_825.vcd");
  if(my_type==3 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_826.vcd");
  if(my_type==3 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_827.vcd");
  if(my_type==3 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_828.vcd");
  if(my_type==3 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_829.vcd");
  if(my_type==3 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_830.vcd");
  if(my_type==3 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_831.vcd");
  if(my_type==3 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_832.vcd");
  if(my_type==3 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_833.vcd");
  if(my_type==3 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_834.vcd");
  if(my_type==3 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_835.vcd");
  if(my_type==3 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_836.vcd");
  if(my_type==3 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_837.vcd");
  if(my_type==3 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_838.vcd");
  if(my_type==3 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_839.vcd");
  if(my_type==3 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_840.vcd");
  if(my_type==3 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_841.vcd");
  if(my_type==3 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_842.vcd");
  if(my_type==3 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_843.vcd");
  if(my_type==3 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_844.vcd");
  if(my_type==3 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_845.vcd");
  if(my_type==3 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_846.vcd");
  if(my_type==3 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_847.vcd");
  if(my_type==3 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_848.vcd");
  if(my_type==3 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_849.vcd");
  if(my_type==3 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_850.vcd");
  if(my_type==3 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_851.vcd");
  if(my_type==3 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_852.vcd");
  if(my_type==3 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_853.vcd");
  if(my_type==3 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_854.vcd");
  if(my_type==3 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_855.vcd");
  if(my_type==3 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_856.vcd");
  if(my_type==3 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_857.vcd");
  if(my_type==3 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_858.vcd");
  if(my_type==3 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_859.vcd");
  if(my_type==3 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_860.vcd");
  if(my_type==3 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_861.vcd");
  if(my_type==3 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_862.vcd");
  if(my_type==3 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_863.vcd");
  if(my_type==3 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_864.vcd");
  if(my_type==3 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_865.vcd");
  if(my_type==3 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_866.vcd");
  if(my_type==3 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_867.vcd");
  if(my_type==3 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_868.vcd");
  if(my_type==3 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_869.vcd");
  if(my_type==3 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_870.vcd");
  if(my_type==3 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_871.vcd");
  if(my_type==3 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_872.vcd");
  if(my_type==3 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_873.vcd");
  if(my_type==3 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_874.vcd");
  if(my_type==3 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_875.vcd");
  if(my_type==3 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_876.vcd");
  if(my_type==3 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_877.vcd");
  if(my_type==3 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_878.vcd");
  if(my_type==3 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_879.vcd");
  if(my_type==3 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_880.vcd");
  if(my_type==3 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_881.vcd");
  if(my_type==3 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_882.vcd");
  if(my_type==3 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_883.vcd");
  if(my_type==3 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_884.vcd");
  if(my_type==3 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_885.vcd");
  if(my_type==3 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_886.vcd");
  if(my_type==3 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_887.vcd");
  if(my_type==3 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_888.vcd");
  if(my_type==3 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_889.vcd");
  if(my_type==3 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_890.vcd");
  if(my_type==3 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_891.vcd");
  if(my_type==3 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_892.vcd");
  if(my_type==3 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_893.vcd");
  if(my_type==3 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_894.vcd");
  if(my_type==3 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_895.vcd");
  if(my_type==3 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_896.vcd");
  if(my_type==3 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_897.vcd");
  if(my_type==3 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_898.vcd");
  if(my_type==3 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_899.vcd");
  if(my_type==3 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_900.vcd");
  if(my_type==3 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_901.vcd");
  if(my_type==3 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_902.vcd");
  if(my_type==3 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_903.vcd");
  if(my_type==3 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_904.vcd");
  if(my_type==3 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_905.vcd");
  if(my_type==3 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_906.vcd");
  if(my_type==3 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_907.vcd");
  if(my_type==3 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_908.vcd");
  if(my_type==3 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_909.vcd");
  if(my_type==3 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_910.vcd");
  if(my_type==3 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_911.vcd");
  if(my_type==3 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_912.vcd");
  if(my_type==3 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_913.vcd");
  if(my_type==3 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_914.vcd");
  if(my_type==3 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_915.vcd");
  if(my_type==3 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_916.vcd");
  if(my_type==3 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_917.vcd");
  if(my_type==3 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_918.vcd");
  if(my_type==3 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_919.vcd");
  if(my_type==3 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_920.vcd");
  if(my_type==3 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_921.vcd");
  if(my_type==3 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_922.vcd");
  if(my_type==3 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_923.vcd");
  if(my_type==3 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_924.vcd");
  if(my_type==3 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_925.vcd");
  if(my_type==3 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_926.vcd");
  if(my_type==3 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_927.vcd");
  if(my_type==3 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_928.vcd");
  if(my_type==3 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_929.vcd");
  if(my_type==3 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_930.vcd");
  if(my_type==3 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_931.vcd");
  if(my_type==3 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_932.vcd");
  if(my_type==3 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_933.vcd");
  if(my_type==3 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_934.vcd");
  if(my_type==3 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_935.vcd");
  if(my_type==3 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_936.vcd");
  if(my_type==3 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_937.vcd");
  if(my_type==3 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_938.vcd");
  if(my_type==3 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_939.vcd");
  if(my_type==3 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_940.vcd");
  if(my_type==3 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_941.vcd");
  if(my_type==3 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_942.vcd");
  if(my_type==3 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_943.vcd");
  if(my_type==3 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_944.vcd");
  if(my_type==3 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_945.vcd");
  if(my_type==3 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_946.vcd");
  if(my_type==3 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_947.vcd");
  if(my_type==3 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_948.vcd");
  if(my_type==3 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_949.vcd");
  if(my_type==3 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_950.vcd");
  if(my_type==3 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_951.vcd");
  if(my_type==3 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_952.vcd");
  if(my_type==3 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_953.vcd");
  if(my_type==3 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_954.vcd");
  if(my_type==3 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_955.vcd");
  if(my_type==3 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_956.vcd");
  if(my_type==3 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_957.vcd");
  if(my_type==3 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_958.vcd");
  if(my_type==3 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_959.vcd");
  if(my_type==3 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_960.vcd");
  if(my_type==3 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_961.vcd");
  if(my_type==3 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_962.vcd");
  if(my_type==3 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_963.vcd");
  if(my_type==3 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_964.vcd");
  if(my_type==3 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_965.vcd");
  if(my_type==3 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_966.vcd");
  if(my_type==3 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_967.vcd");
  if(my_type==3 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_968.vcd");
  if(my_type==3 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_969.vcd");
  if(my_type==3 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_970.vcd");
  if(my_type==3 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_971.vcd");
  if(my_type==3 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_972.vcd");
  if(my_type==3 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_973.vcd");
  if(my_type==3 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_974.vcd");
  if(my_type==3 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_975.vcd");
  if(my_type==3 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_976.vcd");
  if(my_type==3 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_977.vcd");
  if(my_type==3 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_978.vcd");
  if(my_type==3 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_979.vcd");
  if(my_type==3 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_980.vcd");
  if(my_type==3 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_981.vcd");
  if(my_type==3 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_982.vcd");
  if(my_type==3 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_983.vcd");
  if(my_type==3 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_984.vcd");
  if(my_type==3 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_985.vcd");
  if(my_type==3 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_986.vcd");
  if(my_type==3 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_987.vcd");
  if(my_type==3 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_988.vcd");
  if(my_type==3 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_989.vcd");
  if(my_type==3 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_990.vcd");
  if(my_type==3 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_991.vcd");
  if(my_type==3 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_992.vcd");
  if(my_type==3 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_993.vcd");
  if(my_type==3 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_994.vcd");
  if(my_type==3 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_995.vcd");
  if(my_type==3 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_996.vcd");
  if(my_type==3 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_997.vcd");
  if(my_type==3 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_998.vcd");
  if(my_type==3 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_3_999.vcd");
  if(my_type==4 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_0.vcd");
  if(my_type==4 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_1.vcd");
  if(my_type==4 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_2.vcd");
  if(my_type==4 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_3.vcd");
  if(my_type==4 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_4.vcd");
  if(my_type==4 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_5.vcd");
  if(my_type==4 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_6.vcd");
  if(my_type==4 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_7.vcd");
  if(my_type==4 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_8.vcd");
  if(my_type==4 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_9.vcd");
  if(my_type==4 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_10.vcd");
  if(my_type==4 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_11.vcd");
  if(my_type==4 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_12.vcd");
  if(my_type==4 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_13.vcd");
  if(my_type==4 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_14.vcd");
  if(my_type==4 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_15.vcd");
  if(my_type==4 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_16.vcd");
  if(my_type==4 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_17.vcd");
  if(my_type==4 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_18.vcd");
  if(my_type==4 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_19.vcd");
  if(my_type==4 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_20.vcd");
  if(my_type==4 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_21.vcd");
  if(my_type==4 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_22.vcd");
  if(my_type==4 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_23.vcd");
  if(my_type==4 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_24.vcd");
  if(my_type==4 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_25.vcd");
  if(my_type==4 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_26.vcd");
  if(my_type==4 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_27.vcd");
  if(my_type==4 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_28.vcd");
  if(my_type==4 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_29.vcd");
  if(my_type==4 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_30.vcd");
  if(my_type==4 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_31.vcd");
  if(my_type==4 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_32.vcd");
  if(my_type==4 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_33.vcd");
  if(my_type==4 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_34.vcd");
  if(my_type==4 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_35.vcd");
  if(my_type==4 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_36.vcd");
  if(my_type==4 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_37.vcd");
  if(my_type==4 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_38.vcd");
  if(my_type==4 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_39.vcd");
  if(my_type==4 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_40.vcd");
  if(my_type==4 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_41.vcd");
  if(my_type==4 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_42.vcd");
  if(my_type==4 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_43.vcd");
  if(my_type==4 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_44.vcd");
  if(my_type==4 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_45.vcd");
  if(my_type==4 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_46.vcd");
  if(my_type==4 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_47.vcd");
  if(my_type==4 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_48.vcd");
  if(my_type==4 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_49.vcd");
  if(my_type==4 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_50.vcd");
  if(my_type==4 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_51.vcd");
  if(my_type==4 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_52.vcd");
  if(my_type==4 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_53.vcd");
  if(my_type==4 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_54.vcd");
  if(my_type==4 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_55.vcd");
  if(my_type==4 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_56.vcd");
  if(my_type==4 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_57.vcd");
  if(my_type==4 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_58.vcd");
  if(my_type==4 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_59.vcd");
  if(my_type==4 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_60.vcd");
  if(my_type==4 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_61.vcd");
  if(my_type==4 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_62.vcd");
  if(my_type==4 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_63.vcd");
  if(my_type==4 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_64.vcd");
  if(my_type==4 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_65.vcd");
  if(my_type==4 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_66.vcd");
  if(my_type==4 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_67.vcd");
  if(my_type==4 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_68.vcd");
  if(my_type==4 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_69.vcd");
  if(my_type==4 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_70.vcd");
  if(my_type==4 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_71.vcd");
  if(my_type==4 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_72.vcd");
  if(my_type==4 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_73.vcd");
  if(my_type==4 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_74.vcd");
  if(my_type==4 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_75.vcd");
  if(my_type==4 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_76.vcd");
  if(my_type==4 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_77.vcd");
  if(my_type==4 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_78.vcd");
  if(my_type==4 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_79.vcd");
  if(my_type==4 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_80.vcd");
  if(my_type==4 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_81.vcd");
  if(my_type==4 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_82.vcd");
  if(my_type==4 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_83.vcd");
  if(my_type==4 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_84.vcd");
  if(my_type==4 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_85.vcd");
  if(my_type==4 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_86.vcd");
  if(my_type==4 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_87.vcd");
  if(my_type==4 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_88.vcd");
  if(my_type==4 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_89.vcd");
  if(my_type==4 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_90.vcd");
  if(my_type==4 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_91.vcd");
  if(my_type==4 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_92.vcd");
  if(my_type==4 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_93.vcd");
  if(my_type==4 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_94.vcd");
  if(my_type==4 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_95.vcd");
  if(my_type==4 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_96.vcd");
  if(my_type==4 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_97.vcd");
  if(my_type==4 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_98.vcd");
  if(my_type==4 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_99.vcd");
  if(my_type==4 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_100.vcd");
  if(my_type==4 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_101.vcd");
  if(my_type==4 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_102.vcd");
  if(my_type==4 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_103.vcd");
  if(my_type==4 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_104.vcd");
  if(my_type==4 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_105.vcd");
  if(my_type==4 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_106.vcd");
  if(my_type==4 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_107.vcd");
  if(my_type==4 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_108.vcd");
  if(my_type==4 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_109.vcd");
  if(my_type==4 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_110.vcd");
  if(my_type==4 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_111.vcd");
  if(my_type==4 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_112.vcd");
  if(my_type==4 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_113.vcd");
  if(my_type==4 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_114.vcd");
  if(my_type==4 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_115.vcd");
  if(my_type==4 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_116.vcd");
  if(my_type==4 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_117.vcd");
  if(my_type==4 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_118.vcd");
  if(my_type==4 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_119.vcd");
  if(my_type==4 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_120.vcd");
  if(my_type==4 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_121.vcd");
  if(my_type==4 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_122.vcd");
  if(my_type==4 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_123.vcd");
  if(my_type==4 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_124.vcd");
  if(my_type==4 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_125.vcd");
  if(my_type==4 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_126.vcd");
  if(my_type==4 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_127.vcd");
  if(my_type==4 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_128.vcd");
  if(my_type==4 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_129.vcd");
  if(my_type==4 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_130.vcd");
  if(my_type==4 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_131.vcd");
  if(my_type==4 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_132.vcd");
  if(my_type==4 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_133.vcd");
  if(my_type==4 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_134.vcd");
  if(my_type==4 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_135.vcd");
  if(my_type==4 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_136.vcd");
  if(my_type==4 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_137.vcd");
  if(my_type==4 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_138.vcd");
  if(my_type==4 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_139.vcd");
  if(my_type==4 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_140.vcd");
  if(my_type==4 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_141.vcd");
  if(my_type==4 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_142.vcd");
  if(my_type==4 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_143.vcd");
  if(my_type==4 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_144.vcd");
  if(my_type==4 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_145.vcd");
  if(my_type==4 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_146.vcd");
  if(my_type==4 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_147.vcd");
  if(my_type==4 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_148.vcd");
  if(my_type==4 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_149.vcd");
  if(my_type==4 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_150.vcd");
  if(my_type==4 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_151.vcd");
  if(my_type==4 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_152.vcd");
  if(my_type==4 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_153.vcd");
  if(my_type==4 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_154.vcd");
  if(my_type==4 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_155.vcd");
  if(my_type==4 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_156.vcd");
  if(my_type==4 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_157.vcd");
  if(my_type==4 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_158.vcd");
  if(my_type==4 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_159.vcd");
  if(my_type==4 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_160.vcd");
  if(my_type==4 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_161.vcd");
  if(my_type==4 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_162.vcd");
  if(my_type==4 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_163.vcd");
  if(my_type==4 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_164.vcd");
  if(my_type==4 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_165.vcd");
  if(my_type==4 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_166.vcd");
  if(my_type==4 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_167.vcd");
  if(my_type==4 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_168.vcd");
  if(my_type==4 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_169.vcd");
  if(my_type==4 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_170.vcd");
  if(my_type==4 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_171.vcd");
  if(my_type==4 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_172.vcd");
  if(my_type==4 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_173.vcd");
  if(my_type==4 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_174.vcd");
  if(my_type==4 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_175.vcd");
  if(my_type==4 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_176.vcd");
  if(my_type==4 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_177.vcd");
  if(my_type==4 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_178.vcd");
  if(my_type==4 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_179.vcd");
  if(my_type==4 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_180.vcd");
  if(my_type==4 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_181.vcd");
  if(my_type==4 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_182.vcd");
  if(my_type==4 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_183.vcd");
  if(my_type==4 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_184.vcd");
  if(my_type==4 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_185.vcd");
  if(my_type==4 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_186.vcd");
  if(my_type==4 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_187.vcd");
  if(my_type==4 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_188.vcd");
  if(my_type==4 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_189.vcd");
  if(my_type==4 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_190.vcd");
  if(my_type==4 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_191.vcd");
  if(my_type==4 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_192.vcd");
  if(my_type==4 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_193.vcd");
  if(my_type==4 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_194.vcd");
  if(my_type==4 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_195.vcd");
  if(my_type==4 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_196.vcd");
  if(my_type==4 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_197.vcd");
  if(my_type==4 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_198.vcd");
  if(my_type==4 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_199.vcd");
  if(my_type==4 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_200.vcd");
  if(my_type==4 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_201.vcd");
  if(my_type==4 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_202.vcd");
  if(my_type==4 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_203.vcd");
  if(my_type==4 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_204.vcd");
  if(my_type==4 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_205.vcd");
  if(my_type==4 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_206.vcd");
  if(my_type==4 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_207.vcd");
  if(my_type==4 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_208.vcd");
  if(my_type==4 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_209.vcd");
  if(my_type==4 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_210.vcd");
  if(my_type==4 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_211.vcd");
  if(my_type==4 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_212.vcd");
  if(my_type==4 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_213.vcd");
  if(my_type==4 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_214.vcd");
  if(my_type==4 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_215.vcd");
  if(my_type==4 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_216.vcd");
  if(my_type==4 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_217.vcd");
  if(my_type==4 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_218.vcd");
  if(my_type==4 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_219.vcd");
  if(my_type==4 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_220.vcd");
  if(my_type==4 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_221.vcd");
  if(my_type==4 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_222.vcd");
  if(my_type==4 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_223.vcd");
  if(my_type==4 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_224.vcd");
  if(my_type==4 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_225.vcd");
  if(my_type==4 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_226.vcd");
  if(my_type==4 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_227.vcd");
  if(my_type==4 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_228.vcd");
  if(my_type==4 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_229.vcd");
  if(my_type==4 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_230.vcd");
  if(my_type==4 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_231.vcd");
  if(my_type==4 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_232.vcd");
  if(my_type==4 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_233.vcd");
  if(my_type==4 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_234.vcd");
  if(my_type==4 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_235.vcd");
  if(my_type==4 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_236.vcd");
  if(my_type==4 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_237.vcd");
  if(my_type==4 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_238.vcd");
  if(my_type==4 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_239.vcd");
  if(my_type==4 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_240.vcd");
  if(my_type==4 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_241.vcd");
  if(my_type==4 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_242.vcd");
  if(my_type==4 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_243.vcd");
  if(my_type==4 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_244.vcd");
  if(my_type==4 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_245.vcd");
  if(my_type==4 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_246.vcd");
  if(my_type==4 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_247.vcd");
  if(my_type==4 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_248.vcd");
  if(my_type==4 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_249.vcd");
  if(my_type==4 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_250.vcd");
  if(my_type==4 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_251.vcd");
  if(my_type==4 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_252.vcd");
  if(my_type==4 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_253.vcd");
  if(my_type==4 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_254.vcd");
  if(my_type==4 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_255.vcd");
  if(my_type==4 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_256.vcd");
  if(my_type==4 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_257.vcd");
  if(my_type==4 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_258.vcd");
  if(my_type==4 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_259.vcd");
  if(my_type==4 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_260.vcd");
  if(my_type==4 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_261.vcd");
  if(my_type==4 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_262.vcd");
  if(my_type==4 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_263.vcd");
  if(my_type==4 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_264.vcd");
  if(my_type==4 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_265.vcd");
  if(my_type==4 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_266.vcd");
  if(my_type==4 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_267.vcd");
  if(my_type==4 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_268.vcd");
  if(my_type==4 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_269.vcd");
  if(my_type==4 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_270.vcd");
  if(my_type==4 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_271.vcd");
  if(my_type==4 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_272.vcd");
  if(my_type==4 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_273.vcd");
  if(my_type==4 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_274.vcd");
  if(my_type==4 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_275.vcd");
  if(my_type==4 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_276.vcd");
  if(my_type==4 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_277.vcd");
  if(my_type==4 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_278.vcd");
  if(my_type==4 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_279.vcd");
  if(my_type==4 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_280.vcd");
  if(my_type==4 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_281.vcd");
  if(my_type==4 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_282.vcd");
  if(my_type==4 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_283.vcd");
  if(my_type==4 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_284.vcd");
  if(my_type==4 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_285.vcd");
  if(my_type==4 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_286.vcd");
  if(my_type==4 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_287.vcd");
  if(my_type==4 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_288.vcd");
  if(my_type==4 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_289.vcd");
  if(my_type==4 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_290.vcd");
  if(my_type==4 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_291.vcd");
  if(my_type==4 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_292.vcd");
  if(my_type==4 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_293.vcd");
  if(my_type==4 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_294.vcd");
  if(my_type==4 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_295.vcd");
  if(my_type==4 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_296.vcd");
  if(my_type==4 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_297.vcd");
  if(my_type==4 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_298.vcd");
  if(my_type==4 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_299.vcd");
  if(my_type==4 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_300.vcd");
  if(my_type==4 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_301.vcd");
  if(my_type==4 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_302.vcd");
  if(my_type==4 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_303.vcd");
  if(my_type==4 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_304.vcd");
  if(my_type==4 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_305.vcd");
  if(my_type==4 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_306.vcd");
  if(my_type==4 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_307.vcd");
  if(my_type==4 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_308.vcd");
  if(my_type==4 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_309.vcd");
  if(my_type==4 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_310.vcd");
  if(my_type==4 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_311.vcd");
  if(my_type==4 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_312.vcd");
  if(my_type==4 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_313.vcd");
  if(my_type==4 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_314.vcd");
  if(my_type==4 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_315.vcd");
  if(my_type==4 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_316.vcd");
  if(my_type==4 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_317.vcd");
  if(my_type==4 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_318.vcd");
  if(my_type==4 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_319.vcd");
  if(my_type==4 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_320.vcd");
  if(my_type==4 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_321.vcd");
  if(my_type==4 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_322.vcd");
  if(my_type==4 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_323.vcd");
  if(my_type==4 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_324.vcd");
  if(my_type==4 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_325.vcd");
  if(my_type==4 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_326.vcd");
  if(my_type==4 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_327.vcd");
  if(my_type==4 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_328.vcd");
  if(my_type==4 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_329.vcd");
  if(my_type==4 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_330.vcd");
  if(my_type==4 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_331.vcd");
  if(my_type==4 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_332.vcd");
  if(my_type==4 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_333.vcd");
  if(my_type==4 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_334.vcd");
  if(my_type==4 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_335.vcd");
  if(my_type==4 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_336.vcd");
  if(my_type==4 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_337.vcd");
  if(my_type==4 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_338.vcd");
  if(my_type==4 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_339.vcd");
  if(my_type==4 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_340.vcd");
  if(my_type==4 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_341.vcd");
  if(my_type==4 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_342.vcd");
  if(my_type==4 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_343.vcd");
  if(my_type==4 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_344.vcd");
  if(my_type==4 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_345.vcd");
  if(my_type==4 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_346.vcd");
  if(my_type==4 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_347.vcd");
  if(my_type==4 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_348.vcd");
  if(my_type==4 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_349.vcd");
  if(my_type==4 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_350.vcd");
  if(my_type==4 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_351.vcd");
  if(my_type==4 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_352.vcd");
  if(my_type==4 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_353.vcd");
  if(my_type==4 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_354.vcd");
  if(my_type==4 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_355.vcd");
  if(my_type==4 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_356.vcd");
  if(my_type==4 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_357.vcd");
  if(my_type==4 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_358.vcd");
  if(my_type==4 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_359.vcd");
  if(my_type==4 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_360.vcd");
  if(my_type==4 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_361.vcd");
  if(my_type==4 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_362.vcd");
  if(my_type==4 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_363.vcd");
  if(my_type==4 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_364.vcd");
  if(my_type==4 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_365.vcd");
  if(my_type==4 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_366.vcd");
  if(my_type==4 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_367.vcd");
  if(my_type==4 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_368.vcd");
  if(my_type==4 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_369.vcd");
  if(my_type==4 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_370.vcd");
  if(my_type==4 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_371.vcd");
  if(my_type==4 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_372.vcd");
  if(my_type==4 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_373.vcd");
  if(my_type==4 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_374.vcd");
  if(my_type==4 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_375.vcd");
  if(my_type==4 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_376.vcd");
  if(my_type==4 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_377.vcd");
  if(my_type==4 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_378.vcd");
  if(my_type==4 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_379.vcd");
  if(my_type==4 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_380.vcd");
  if(my_type==4 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_381.vcd");
  if(my_type==4 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_382.vcd");
  if(my_type==4 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_383.vcd");
  if(my_type==4 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_384.vcd");
  if(my_type==4 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_385.vcd");
  if(my_type==4 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_386.vcd");
  if(my_type==4 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_387.vcd");
  if(my_type==4 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_388.vcd");
  if(my_type==4 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_389.vcd");
  if(my_type==4 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_390.vcd");
  if(my_type==4 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_391.vcd");
  if(my_type==4 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_392.vcd");
  if(my_type==4 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_393.vcd");
  if(my_type==4 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_394.vcd");
  if(my_type==4 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_395.vcd");
  if(my_type==4 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_396.vcd");
  if(my_type==4 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_397.vcd");
  if(my_type==4 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_398.vcd");
  if(my_type==4 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_399.vcd");
  if(my_type==4 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_400.vcd");
  if(my_type==4 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_401.vcd");
  if(my_type==4 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_402.vcd");
  if(my_type==4 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_403.vcd");
  if(my_type==4 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_404.vcd");
  if(my_type==4 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_405.vcd");
  if(my_type==4 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_406.vcd");
  if(my_type==4 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_407.vcd");
  if(my_type==4 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_408.vcd");
  if(my_type==4 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_409.vcd");
  if(my_type==4 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_410.vcd");
  if(my_type==4 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_411.vcd");
  if(my_type==4 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_412.vcd");
  if(my_type==4 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_413.vcd");
  if(my_type==4 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_414.vcd");
  if(my_type==4 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_415.vcd");
  if(my_type==4 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_416.vcd");
  if(my_type==4 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_417.vcd");
  if(my_type==4 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_418.vcd");
  if(my_type==4 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_419.vcd");
  if(my_type==4 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_420.vcd");
  if(my_type==4 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_421.vcd");
  if(my_type==4 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_422.vcd");
  if(my_type==4 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_423.vcd");
  if(my_type==4 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_424.vcd");
  if(my_type==4 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_425.vcd");
  if(my_type==4 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_426.vcd");
  if(my_type==4 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_427.vcd");
  if(my_type==4 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_428.vcd");
  if(my_type==4 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_429.vcd");
  if(my_type==4 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_430.vcd");
  if(my_type==4 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_431.vcd");
  if(my_type==4 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_432.vcd");
  if(my_type==4 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_433.vcd");
  if(my_type==4 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_434.vcd");
  if(my_type==4 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_435.vcd");
  if(my_type==4 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_436.vcd");
  if(my_type==4 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_437.vcd");
  if(my_type==4 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_438.vcd");
  if(my_type==4 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_439.vcd");
  if(my_type==4 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_440.vcd");
  if(my_type==4 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_441.vcd");
  if(my_type==4 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_442.vcd");
  if(my_type==4 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_443.vcd");
  if(my_type==4 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_444.vcd");
  if(my_type==4 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_445.vcd");
  if(my_type==4 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_446.vcd");
  if(my_type==4 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_447.vcd");
  if(my_type==4 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_448.vcd");
  if(my_type==4 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_449.vcd");
  if(my_type==4 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_450.vcd");
  if(my_type==4 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_451.vcd");
  if(my_type==4 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_452.vcd");
  if(my_type==4 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_453.vcd");
  if(my_type==4 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_454.vcd");
  if(my_type==4 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_455.vcd");
  if(my_type==4 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_456.vcd");
  if(my_type==4 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_457.vcd");
  if(my_type==4 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_458.vcd");
  if(my_type==4 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_459.vcd");
  if(my_type==4 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_460.vcd");
  if(my_type==4 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_461.vcd");
  if(my_type==4 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_462.vcd");
  if(my_type==4 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_463.vcd");
  if(my_type==4 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_464.vcd");
  if(my_type==4 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_465.vcd");
  if(my_type==4 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_466.vcd");
  if(my_type==4 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_467.vcd");
  if(my_type==4 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_468.vcd");
  if(my_type==4 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_469.vcd");
  if(my_type==4 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_470.vcd");
  if(my_type==4 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_471.vcd");
  if(my_type==4 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_472.vcd");
  if(my_type==4 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_473.vcd");
  if(my_type==4 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_474.vcd");
  if(my_type==4 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_475.vcd");
  if(my_type==4 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_476.vcd");
  if(my_type==4 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_477.vcd");
  if(my_type==4 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_478.vcd");
  if(my_type==4 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_479.vcd");
  if(my_type==4 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_480.vcd");
  if(my_type==4 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_481.vcd");
  if(my_type==4 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_482.vcd");
  if(my_type==4 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_483.vcd");
  if(my_type==4 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_484.vcd");
  if(my_type==4 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_485.vcd");
  if(my_type==4 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_486.vcd");
  if(my_type==4 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_487.vcd");
  if(my_type==4 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_488.vcd");
  if(my_type==4 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_489.vcd");
  if(my_type==4 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_490.vcd");
  if(my_type==4 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_491.vcd");
  if(my_type==4 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_492.vcd");
  if(my_type==4 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_493.vcd");
  if(my_type==4 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_494.vcd");
  if(my_type==4 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_495.vcd");
  if(my_type==4 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_496.vcd");
  if(my_type==4 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_497.vcd");
  if(my_type==4 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_498.vcd");
  if(my_type==4 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_499.vcd");
  if(my_type==4 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_500.vcd");
  if(my_type==4 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_501.vcd");
  if(my_type==4 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_502.vcd");
  if(my_type==4 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_503.vcd");
  if(my_type==4 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_504.vcd");
  if(my_type==4 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_505.vcd");
  if(my_type==4 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_506.vcd");
  if(my_type==4 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_507.vcd");
  if(my_type==4 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_508.vcd");
  if(my_type==4 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_509.vcd");
  if(my_type==4 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_510.vcd");
  if(my_type==4 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_511.vcd");
  if(my_type==4 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_512.vcd");
  if(my_type==4 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_513.vcd");
  if(my_type==4 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_514.vcd");
  if(my_type==4 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_515.vcd");
  if(my_type==4 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_516.vcd");
  if(my_type==4 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_517.vcd");
  if(my_type==4 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_518.vcd");
  if(my_type==4 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_519.vcd");
  if(my_type==4 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_520.vcd");
  if(my_type==4 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_521.vcd");
  if(my_type==4 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_522.vcd");
  if(my_type==4 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_523.vcd");
  if(my_type==4 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_524.vcd");
  if(my_type==4 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_525.vcd");
  if(my_type==4 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_526.vcd");
  if(my_type==4 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_527.vcd");
  if(my_type==4 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_528.vcd");
  if(my_type==4 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_529.vcd");
  if(my_type==4 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_530.vcd");
  if(my_type==4 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_531.vcd");
  if(my_type==4 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_532.vcd");
  if(my_type==4 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_533.vcd");
  if(my_type==4 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_534.vcd");
  if(my_type==4 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_535.vcd");
  if(my_type==4 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_536.vcd");
  if(my_type==4 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_537.vcd");
  if(my_type==4 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_538.vcd");
  if(my_type==4 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_539.vcd");
  if(my_type==4 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_540.vcd");
  if(my_type==4 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_541.vcd");
  if(my_type==4 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_542.vcd");
  if(my_type==4 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_543.vcd");
  if(my_type==4 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_544.vcd");
  if(my_type==4 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_545.vcd");
  if(my_type==4 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_546.vcd");
  if(my_type==4 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_547.vcd");
  if(my_type==4 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_548.vcd");
  if(my_type==4 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_549.vcd");
  if(my_type==4 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_550.vcd");
  if(my_type==4 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_551.vcd");
  if(my_type==4 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_552.vcd");
  if(my_type==4 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_553.vcd");
  if(my_type==4 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_554.vcd");
  if(my_type==4 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_555.vcd");
  if(my_type==4 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_556.vcd");
  if(my_type==4 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_557.vcd");
  if(my_type==4 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_558.vcd");
  if(my_type==4 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_559.vcd");
  if(my_type==4 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_560.vcd");
  if(my_type==4 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_561.vcd");
  if(my_type==4 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_562.vcd");
  if(my_type==4 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_563.vcd");
  if(my_type==4 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_564.vcd");
  if(my_type==4 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_565.vcd");
  if(my_type==4 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_566.vcd");
  if(my_type==4 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_567.vcd");
  if(my_type==4 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_568.vcd");
  if(my_type==4 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_569.vcd");
  if(my_type==4 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_570.vcd");
  if(my_type==4 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_571.vcd");
  if(my_type==4 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_572.vcd");
  if(my_type==4 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_573.vcd");
  if(my_type==4 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_574.vcd");
  if(my_type==4 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_575.vcd");
  if(my_type==4 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_576.vcd");
  if(my_type==4 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_577.vcd");
  if(my_type==4 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_578.vcd");
  if(my_type==4 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_579.vcd");
  if(my_type==4 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_580.vcd");
  if(my_type==4 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_581.vcd");
  if(my_type==4 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_582.vcd");
  if(my_type==4 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_583.vcd");
  if(my_type==4 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_584.vcd");
  if(my_type==4 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_585.vcd");
  if(my_type==4 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_586.vcd");
  if(my_type==4 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_587.vcd");
  if(my_type==4 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_588.vcd");
  if(my_type==4 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_589.vcd");
  if(my_type==4 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_590.vcd");
  if(my_type==4 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_591.vcd");
  if(my_type==4 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_592.vcd");
  if(my_type==4 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_593.vcd");
  if(my_type==4 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_594.vcd");
  if(my_type==4 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_595.vcd");
  if(my_type==4 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_596.vcd");
  if(my_type==4 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_597.vcd");
  if(my_type==4 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_598.vcd");
  if(my_type==4 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_599.vcd");
  if(my_type==4 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_600.vcd");
  if(my_type==4 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_601.vcd");
  if(my_type==4 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_602.vcd");
  if(my_type==4 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_603.vcd");
  if(my_type==4 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_604.vcd");
  if(my_type==4 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_605.vcd");
  if(my_type==4 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_606.vcd");
  if(my_type==4 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_607.vcd");
  if(my_type==4 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_608.vcd");
  if(my_type==4 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_609.vcd");
  if(my_type==4 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_610.vcd");
  if(my_type==4 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_611.vcd");
  if(my_type==4 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_612.vcd");
  if(my_type==4 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_613.vcd");
  if(my_type==4 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_614.vcd");
  if(my_type==4 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_615.vcd");
  if(my_type==4 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_616.vcd");
  if(my_type==4 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_617.vcd");
  if(my_type==4 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_618.vcd");
  if(my_type==4 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_619.vcd");
  if(my_type==4 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_620.vcd");
  if(my_type==4 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_621.vcd");
  if(my_type==4 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_622.vcd");
  if(my_type==4 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_623.vcd");
  if(my_type==4 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_624.vcd");
  if(my_type==4 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_625.vcd");
  if(my_type==4 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_626.vcd");
  if(my_type==4 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_627.vcd");
  if(my_type==4 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_628.vcd");
  if(my_type==4 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_629.vcd");
  if(my_type==4 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_630.vcd");
  if(my_type==4 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_631.vcd");
  if(my_type==4 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_632.vcd");
  if(my_type==4 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_633.vcd");
  if(my_type==4 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_634.vcd");
  if(my_type==4 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_635.vcd");
  if(my_type==4 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_636.vcd");
  if(my_type==4 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_637.vcd");
  if(my_type==4 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_638.vcd");
  if(my_type==4 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_639.vcd");
  if(my_type==4 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_640.vcd");
  if(my_type==4 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_641.vcd");
  if(my_type==4 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_642.vcd");
  if(my_type==4 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_643.vcd");
  if(my_type==4 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_644.vcd");
  if(my_type==4 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_645.vcd");
  if(my_type==4 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_646.vcd");
  if(my_type==4 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_647.vcd");
  if(my_type==4 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_648.vcd");
  if(my_type==4 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_649.vcd");
  if(my_type==4 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_650.vcd");
  if(my_type==4 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_651.vcd");
  if(my_type==4 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_652.vcd");
  if(my_type==4 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_653.vcd");
  if(my_type==4 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_654.vcd");
  if(my_type==4 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_655.vcd");
  if(my_type==4 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_656.vcd");
  if(my_type==4 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_657.vcd");
  if(my_type==4 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_658.vcd");
  if(my_type==4 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_659.vcd");
  if(my_type==4 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_660.vcd");
  if(my_type==4 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_661.vcd");
  if(my_type==4 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_662.vcd");
  if(my_type==4 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_663.vcd");
  if(my_type==4 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_664.vcd");
  if(my_type==4 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_665.vcd");
  if(my_type==4 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_666.vcd");
  if(my_type==4 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_667.vcd");
  if(my_type==4 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_668.vcd");
  if(my_type==4 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_669.vcd");
  if(my_type==4 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_670.vcd");
  if(my_type==4 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_671.vcd");
  if(my_type==4 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_672.vcd");
  if(my_type==4 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_673.vcd");
  if(my_type==4 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_674.vcd");
  if(my_type==4 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_675.vcd");
  if(my_type==4 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_676.vcd");
  if(my_type==4 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_677.vcd");
  if(my_type==4 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_678.vcd");
  if(my_type==4 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_679.vcd");
  if(my_type==4 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_680.vcd");
  if(my_type==4 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_681.vcd");
  if(my_type==4 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_682.vcd");
  if(my_type==4 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_683.vcd");
  if(my_type==4 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_684.vcd");
  if(my_type==4 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_685.vcd");
  if(my_type==4 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_686.vcd");
  if(my_type==4 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_687.vcd");
  if(my_type==4 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_688.vcd");
  if(my_type==4 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_689.vcd");
  if(my_type==4 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_690.vcd");
  if(my_type==4 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_691.vcd");
  if(my_type==4 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_692.vcd");
  if(my_type==4 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_693.vcd");
  if(my_type==4 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_694.vcd");
  if(my_type==4 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_695.vcd");
  if(my_type==4 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_696.vcd");
  if(my_type==4 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_697.vcd");
  if(my_type==4 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_698.vcd");
  if(my_type==4 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_699.vcd");
  if(my_type==4 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_700.vcd");
  if(my_type==4 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_701.vcd");
  if(my_type==4 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_702.vcd");
  if(my_type==4 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_703.vcd");
  if(my_type==4 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_704.vcd");
  if(my_type==4 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_705.vcd");
  if(my_type==4 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_706.vcd");
  if(my_type==4 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_707.vcd");
  if(my_type==4 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_708.vcd");
  if(my_type==4 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_709.vcd");
  if(my_type==4 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_710.vcd");
  if(my_type==4 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_711.vcd");
  if(my_type==4 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_712.vcd");
  if(my_type==4 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_713.vcd");
  if(my_type==4 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_714.vcd");
  if(my_type==4 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_715.vcd");
  if(my_type==4 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_716.vcd");
  if(my_type==4 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_717.vcd");
  if(my_type==4 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_718.vcd");
  if(my_type==4 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_719.vcd");
  if(my_type==4 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_720.vcd");
  if(my_type==4 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_721.vcd");
  if(my_type==4 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_722.vcd");
  if(my_type==4 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_723.vcd");
  if(my_type==4 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_724.vcd");
  if(my_type==4 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_725.vcd");
  if(my_type==4 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_726.vcd");
  if(my_type==4 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_727.vcd");
  if(my_type==4 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_728.vcd");
  if(my_type==4 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_729.vcd");
  if(my_type==4 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_730.vcd");
  if(my_type==4 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_731.vcd");
  if(my_type==4 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_732.vcd");
  if(my_type==4 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_733.vcd");
  if(my_type==4 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_734.vcd");
  if(my_type==4 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_735.vcd");
  if(my_type==4 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_736.vcd");
  if(my_type==4 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_737.vcd");
  if(my_type==4 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_738.vcd");
  if(my_type==4 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_739.vcd");
  if(my_type==4 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_740.vcd");
  if(my_type==4 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_741.vcd");
  if(my_type==4 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_742.vcd");
  if(my_type==4 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_743.vcd");
  if(my_type==4 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_744.vcd");
  if(my_type==4 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_745.vcd");
  if(my_type==4 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_746.vcd");
  if(my_type==4 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_747.vcd");
  if(my_type==4 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_748.vcd");
  if(my_type==4 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_749.vcd");
  if(my_type==4 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_750.vcd");
  if(my_type==4 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_751.vcd");
  if(my_type==4 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_752.vcd");
  if(my_type==4 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_753.vcd");
  if(my_type==4 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_754.vcd");
  if(my_type==4 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_755.vcd");
  if(my_type==4 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_756.vcd");
  if(my_type==4 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_757.vcd");
  if(my_type==4 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_758.vcd");
  if(my_type==4 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_759.vcd");
  if(my_type==4 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_760.vcd");
  if(my_type==4 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_761.vcd");
  if(my_type==4 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_762.vcd");
  if(my_type==4 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_763.vcd");
  if(my_type==4 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_764.vcd");
  if(my_type==4 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_765.vcd");
  if(my_type==4 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_766.vcd");
  if(my_type==4 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_767.vcd");
  if(my_type==4 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_768.vcd");
  if(my_type==4 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_769.vcd");
  if(my_type==4 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_770.vcd");
  if(my_type==4 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_771.vcd");
  if(my_type==4 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_772.vcd");
  if(my_type==4 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_773.vcd");
  if(my_type==4 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_774.vcd");
  if(my_type==4 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_775.vcd");
  if(my_type==4 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_776.vcd");
  if(my_type==4 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_777.vcd");
  if(my_type==4 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_778.vcd");
  if(my_type==4 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_779.vcd");
  if(my_type==4 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_780.vcd");
  if(my_type==4 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_781.vcd");
  if(my_type==4 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_782.vcd");
  if(my_type==4 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_783.vcd");
  if(my_type==4 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_784.vcd");
  if(my_type==4 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_785.vcd");
  if(my_type==4 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_786.vcd");
  if(my_type==4 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_787.vcd");
  if(my_type==4 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_788.vcd");
  if(my_type==4 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_789.vcd");
  if(my_type==4 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_790.vcd");
  if(my_type==4 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_791.vcd");
  if(my_type==4 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_792.vcd");
  if(my_type==4 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_793.vcd");
  if(my_type==4 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_794.vcd");
  if(my_type==4 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_795.vcd");
  if(my_type==4 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_796.vcd");
  if(my_type==4 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_797.vcd");
  if(my_type==4 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_798.vcd");
  if(my_type==4 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_799.vcd");
  if(my_type==4 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_800.vcd");
  if(my_type==4 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_801.vcd");
  if(my_type==4 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_802.vcd");
  if(my_type==4 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_803.vcd");
  if(my_type==4 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_804.vcd");
  if(my_type==4 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_805.vcd");
  if(my_type==4 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_806.vcd");
  if(my_type==4 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_807.vcd");
  if(my_type==4 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_808.vcd");
  if(my_type==4 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_809.vcd");
  if(my_type==4 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_810.vcd");
  if(my_type==4 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_811.vcd");
  if(my_type==4 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_812.vcd");
  if(my_type==4 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_813.vcd");
  if(my_type==4 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_814.vcd");
  if(my_type==4 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_815.vcd");
  if(my_type==4 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_816.vcd");
  if(my_type==4 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_817.vcd");
  if(my_type==4 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_818.vcd");
  if(my_type==4 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_819.vcd");
  if(my_type==4 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_820.vcd");
  if(my_type==4 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_821.vcd");
  if(my_type==4 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_822.vcd");
  if(my_type==4 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_823.vcd");
  if(my_type==4 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_824.vcd");
  if(my_type==4 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_825.vcd");
  if(my_type==4 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_826.vcd");
  if(my_type==4 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_827.vcd");
  if(my_type==4 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_828.vcd");
  if(my_type==4 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_829.vcd");
  if(my_type==4 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_830.vcd");
  if(my_type==4 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_831.vcd");
  if(my_type==4 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_832.vcd");
  if(my_type==4 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_833.vcd");
  if(my_type==4 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_834.vcd");
  if(my_type==4 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_835.vcd");
  if(my_type==4 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_836.vcd");
  if(my_type==4 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_837.vcd");
  if(my_type==4 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_838.vcd");
  if(my_type==4 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_839.vcd");
  if(my_type==4 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_840.vcd");
  if(my_type==4 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_841.vcd");
  if(my_type==4 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_842.vcd");
  if(my_type==4 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_843.vcd");
  if(my_type==4 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_844.vcd");
  if(my_type==4 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_845.vcd");
  if(my_type==4 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_846.vcd");
  if(my_type==4 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_847.vcd");
  if(my_type==4 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_848.vcd");
  if(my_type==4 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_849.vcd");
  if(my_type==4 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_850.vcd");
  if(my_type==4 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_851.vcd");
  if(my_type==4 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_852.vcd");
  if(my_type==4 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_853.vcd");
  if(my_type==4 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_854.vcd");
  if(my_type==4 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_855.vcd");
  if(my_type==4 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_856.vcd");
  if(my_type==4 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_857.vcd");
  if(my_type==4 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_858.vcd");
  if(my_type==4 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_859.vcd");
  if(my_type==4 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_860.vcd");
  if(my_type==4 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_861.vcd");
  if(my_type==4 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_862.vcd");
  if(my_type==4 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_863.vcd");
  if(my_type==4 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_864.vcd");
  if(my_type==4 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_865.vcd");
  if(my_type==4 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_866.vcd");
  if(my_type==4 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_867.vcd");
  if(my_type==4 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_868.vcd");
  if(my_type==4 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_869.vcd");
  if(my_type==4 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_870.vcd");
  if(my_type==4 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_871.vcd");
  if(my_type==4 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_872.vcd");
  if(my_type==4 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_873.vcd");
  if(my_type==4 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_874.vcd");
  if(my_type==4 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_875.vcd");
  if(my_type==4 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_876.vcd");
  if(my_type==4 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_877.vcd");
  if(my_type==4 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_878.vcd");
  if(my_type==4 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_879.vcd");
  if(my_type==4 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_880.vcd");
  if(my_type==4 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_881.vcd");
  if(my_type==4 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_882.vcd");
  if(my_type==4 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_883.vcd");
  if(my_type==4 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_884.vcd");
  if(my_type==4 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_885.vcd");
  if(my_type==4 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_886.vcd");
  if(my_type==4 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_887.vcd");
  if(my_type==4 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_888.vcd");
  if(my_type==4 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_889.vcd");
  if(my_type==4 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_890.vcd");
  if(my_type==4 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_891.vcd");
  if(my_type==4 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_892.vcd");
  if(my_type==4 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_893.vcd");
  if(my_type==4 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_894.vcd");
  if(my_type==4 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_895.vcd");
  if(my_type==4 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_896.vcd");
  if(my_type==4 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_897.vcd");
  if(my_type==4 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_898.vcd");
  if(my_type==4 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_899.vcd");
  if(my_type==4 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_900.vcd");
  if(my_type==4 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_901.vcd");
  if(my_type==4 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_902.vcd");
  if(my_type==4 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_903.vcd");
  if(my_type==4 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_904.vcd");
  if(my_type==4 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_905.vcd");
  if(my_type==4 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_906.vcd");
  if(my_type==4 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_907.vcd");
  if(my_type==4 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_908.vcd");
  if(my_type==4 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_909.vcd");
  if(my_type==4 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_910.vcd");
  if(my_type==4 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_911.vcd");
  if(my_type==4 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_912.vcd");
  if(my_type==4 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_913.vcd");
  if(my_type==4 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_914.vcd");
  if(my_type==4 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_915.vcd");
  if(my_type==4 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_916.vcd");
  if(my_type==4 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_917.vcd");
  if(my_type==4 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_918.vcd");
  if(my_type==4 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_919.vcd");
  if(my_type==4 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_920.vcd");
  if(my_type==4 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_921.vcd");
  if(my_type==4 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_922.vcd");
  if(my_type==4 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_923.vcd");
  if(my_type==4 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_924.vcd");
  if(my_type==4 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_925.vcd");
  if(my_type==4 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_926.vcd");
  if(my_type==4 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_927.vcd");
  if(my_type==4 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_928.vcd");
  if(my_type==4 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_929.vcd");
  if(my_type==4 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_930.vcd");
  if(my_type==4 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_931.vcd");
  if(my_type==4 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_932.vcd");
  if(my_type==4 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_933.vcd");
  if(my_type==4 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_934.vcd");
  if(my_type==4 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_935.vcd");
  if(my_type==4 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_936.vcd");
  if(my_type==4 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_937.vcd");
  if(my_type==4 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_938.vcd");
  if(my_type==4 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_939.vcd");
  if(my_type==4 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_940.vcd");
  if(my_type==4 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_941.vcd");
  if(my_type==4 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_942.vcd");
  if(my_type==4 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_943.vcd");
  if(my_type==4 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_944.vcd");
  if(my_type==4 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_945.vcd");
  if(my_type==4 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_946.vcd");
  if(my_type==4 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_947.vcd");
  if(my_type==4 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_948.vcd");
  if(my_type==4 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_949.vcd");
  if(my_type==4 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_950.vcd");
  if(my_type==4 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_951.vcd");
  if(my_type==4 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_952.vcd");
  if(my_type==4 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_953.vcd");
  if(my_type==4 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_954.vcd");
  if(my_type==4 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_955.vcd");
  if(my_type==4 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_956.vcd");
  if(my_type==4 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_957.vcd");
  if(my_type==4 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_958.vcd");
  if(my_type==4 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_959.vcd");
  if(my_type==4 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_960.vcd");
  if(my_type==4 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_961.vcd");
  if(my_type==4 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_962.vcd");
  if(my_type==4 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_963.vcd");
  if(my_type==4 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_964.vcd");
  if(my_type==4 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_965.vcd");
  if(my_type==4 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_966.vcd");
  if(my_type==4 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_967.vcd");
  if(my_type==4 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_968.vcd");
  if(my_type==4 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_969.vcd");
  if(my_type==4 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_970.vcd");
  if(my_type==4 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_971.vcd");
  if(my_type==4 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_972.vcd");
  if(my_type==4 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_973.vcd");
  if(my_type==4 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_974.vcd");
  if(my_type==4 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_975.vcd");
  if(my_type==4 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_976.vcd");
  if(my_type==4 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_977.vcd");
  if(my_type==4 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_978.vcd");
  if(my_type==4 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_979.vcd");
  if(my_type==4 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_980.vcd");
  if(my_type==4 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_981.vcd");
  if(my_type==4 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_982.vcd");
  if(my_type==4 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_983.vcd");
  if(my_type==4 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_984.vcd");
  if(my_type==4 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_985.vcd");
  if(my_type==4 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_986.vcd");
  if(my_type==4 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_987.vcd");
  if(my_type==4 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_988.vcd");
  if(my_type==4 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_989.vcd");
  if(my_type==4 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_990.vcd");
  if(my_type==4 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_991.vcd");
  if(my_type==4 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_992.vcd");
  if(my_type==4 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_993.vcd");
  if(my_type==4 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_994.vcd");
  if(my_type==4 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_995.vcd");
  if(my_type==4 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_996.vcd");
  if(my_type==4 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_997.vcd");
  if(my_type==4 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_998.vcd");
  if(my_type==4 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_4_999.vcd");
  if(my_type==5 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_0.vcd");
  if(my_type==5 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_1.vcd");
  if(my_type==5 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_2.vcd");
  if(my_type==5 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_3.vcd");
  if(my_type==5 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_4.vcd");
  if(my_type==5 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_5.vcd");
  if(my_type==5 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_6.vcd");
  if(my_type==5 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_7.vcd");
  if(my_type==5 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_8.vcd");
  if(my_type==5 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_9.vcd");
  if(my_type==5 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_10.vcd");
  if(my_type==5 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_11.vcd");
  if(my_type==5 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_12.vcd");
  if(my_type==5 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_13.vcd");
  if(my_type==5 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_14.vcd");
  if(my_type==5 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_15.vcd");
  if(my_type==5 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_16.vcd");
  if(my_type==5 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_17.vcd");
  if(my_type==5 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_18.vcd");
  if(my_type==5 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_19.vcd");
  if(my_type==5 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_20.vcd");
  if(my_type==5 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_21.vcd");
  if(my_type==5 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_22.vcd");
  if(my_type==5 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_23.vcd");
  if(my_type==5 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_24.vcd");
  if(my_type==5 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_25.vcd");
  if(my_type==5 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_26.vcd");
  if(my_type==5 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_27.vcd");
  if(my_type==5 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_28.vcd");
  if(my_type==5 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_29.vcd");
  if(my_type==5 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_30.vcd");
  if(my_type==5 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_31.vcd");
  if(my_type==5 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_32.vcd");
  if(my_type==5 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_33.vcd");
  if(my_type==5 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_34.vcd");
  if(my_type==5 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_35.vcd");
  if(my_type==5 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_36.vcd");
  if(my_type==5 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_37.vcd");
  if(my_type==5 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_38.vcd");
  if(my_type==5 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_39.vcd");
  if(my_type==5 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_40.vcd");
  if(my_type==5 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_41.vcd");
  if(my_type==5 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_42.vcd");
  if(my_type==5 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_43.vcd");
  if(my_type==5 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_44.vcd");
  if(my_type==5 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_45.vcd");
  if(my_type==5 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_46.vcd");
  if(my_type==5 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_47.vcd");
  if(my_type==5 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_48.vcd");
  if(my_type==5 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_49.vcd");
  if(my_type==5 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_50.vcd");
  if(my_type==5 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_51.vcd");
  if(my_type==5 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_52.vcd");
  if(my_type==5 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_53.vcd");
  if(my_type==5 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_54.vcd");
  if(my_type==5 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_55.vcd");
  if(my_type==5 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_56.vcd");
  if(my_type==5 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_57.vcd");
  if(my_type==5 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_58.vcd");
  if(my_type==5 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_59.vcd");
  if(my_type==5 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_60.vcd");
  if(my_type==5 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_61.vcd");
  if(my_type==5 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_62.vcd");
  if(my_type==5 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_63.vcd");
  if(my_type==5 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_64.vcd");
  if(my_type==5 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_65.vcd");
  if(my_type==5 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_66.vcd");
  if(my_type==5 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_67.vcd");
  if(my_type==5 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_68.vcd");
  if(my_type==5 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_69.vcd");
  if(my_type==5 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_70.vcd");
  if(my_type==5 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_71.vcd");
  if(my_type==5 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_72.vcd");
  if(my_type==5 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_73.vcd");
  if(my_type==5 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_74.vcd");
  if(my_type==5 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_75.vcd");
  if(my_type==5 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_76.vcd");
  if(my_type==5 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_77.vcd");
  if(my_type==5 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_78.vcd");
  if(my_type==5 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_79.vcd");
  if(my_type==5 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_80.vcd");
  if(my_type==5 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_81.vcd");
  if(my_type==5 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_82.vcd");
  if(my_type==5 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_83.vcd");
  if(my_type==5 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_84.vcd");
  if(my_type==5 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_85.vcd");
  if(my_type==5 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_86.vcd");
  if(my_type==5 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_87.vcd");
  if(my_type==5 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_88.vcd");
  if(my_type==5 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_89.vcd");
  if(my_type==5 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_90.vcd");
  if(my_type==5 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_91.vcd");
  if(my_type==5 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_92.vcd");
  if(my_type==5 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_93.vcd");
  if(my_type==5 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_94.vcd");
  if(my_type==5 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_95.vcd");
  if(my_type==5 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_96.vcd");
  if(my_type==5 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_97.vcd");
  if(my_type==5 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_98.vcd");
  if(my_type==5 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_99.vcd");
  if(my_type==5 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_100.vcd");
  if(my_type==5 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_101.vcd");
  if(my_type==5 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_102.vcd");
  if(my_type==5 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_103.vcd");
  if(my_type==5 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_104.vcd");
  if(my_type==5 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_105.vcd");
  if(my_type==5 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_106.vcd");
  if(my_type==5 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_107.vcd");
  if(my_type==5 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_108.vcd");
  if(my_type==5 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_109.vcd");
  if(my_type==5 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_110.vcd");
  if(my_type==5 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_111.vcd");
  if(my_type==5 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_112.vcd");
  if(my_type==5 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_113.vcd");
  if(my_type==5 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_114.vcd");
  if(my_type==5 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_115.vcd");
  if(my_type==5 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_116.vcd");
  if(my_type==5 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_117.vcd");
  if(my_type==5 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_118.vcd");
  if(my_type==5 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_119.vcd");
  if(my_type==5 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_120.vcd");
  if(my_type==5 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_121.vcd");
  if(my_type==5 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_122.vcd");
  if(my_type==5 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_123.vcd");
  if(my_type==5 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_124.vcd");
  if(my_type==5 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_125.vcd");
  if(my_type==5 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_126.vcd");
  if(my_type==5 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_127.vcd");
  if(my_type==5 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_128.vcd");
  if(my_type==5 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_129.vcd");
  if(my_type==5 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_130.vcd");
  if(my_type==5 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_131.vcd");
  if(my_type==5 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_132.vcd");
  if(my_type==5 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_133.vcd");
  if(my_type==5 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_134.vcd");
  if(my_type==5 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_135.vcd");
  if(my_type==5 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_136.vcd");
  if(my_type==5 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_137.vcd");
  if(my_type==5 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_138.vcd");
  if(my_type==5 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_139.vcd");
  if(my_type==5 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_140.vcd");
  if(my_type==5 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_141.vcd");
  if(my_type==5 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_142.vcd");
  if(my_type==5 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_143.vcd");
  if(my_type==5 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_144.vcd");
  if(my_type==5 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_145.vcd");
  if(my_type==5 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_146.vcd");
  if(my_type==5 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_147.vcd");
  if(my_type==5 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_148.vcd");
  if(my_type==5 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_149.vcd");
  if(my_type==5 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_150.vcd");
  if(my_type==5 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_151.vcd");
  if(my_type==5 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_152.vcd");
  if(my_type==5 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_153.vcd");
  if(my_type==5 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_154.vcd");
  if(my_type==5 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_155.vcd");
  if(my_type==5 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_156.vcd");
  if(my_type==5 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_157.vcd");
  if(my_type==5 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_158.vcd");
  if(my_type==5 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_159.vcd");
  if(my_type==5 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_160.vcd");
  if(my_type==5 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_161.vcd");
  if(my_type==5 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_162.vcd");
  if(my_type==5 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_163.vcd");
  if(my_type==5 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_164.vcd");
  if(my_type==5 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_165.vcd");
  if(my_type==5 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_166.vcd");
  if(my_type==5 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_167.vcd");
  if(my_type==5 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_168.vcd");
  if(my_type==5 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_169.vcd");
  if(my_type==5 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_170.vcd");
  if(my_type==5 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_171.vcd");
  if(my_type==5 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_172.vcd");
  if(my_type==5 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_173.vcd");
  if(my_type==5 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_174.vcd");
  if(my_type==5 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_175.vcd");
  if(my_type==5 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_176.vcd");
  if(my_type==5 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_177.vcd");
  if(my_type==5 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_178.vcd");
  if(my_type==5 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_179.vcd");
  if(my_type==5 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_180.vcd");
  if(my_type==5 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_181.vcd");
  if(my_type==5 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_182.vcd");
  if(my_type==5 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_183.vcd");
  if(my_type==5 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_184.vcd");
  if(my_type==5 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_185.vcd");
  if(my_type==5 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_186.vcd");
  if(my_type==5 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_187.vcd");
  if(my_type==5 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_188.vcd");
  if(my_type==5 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_189.vcd");
  if(my_type==5 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_190.vcd");
  if(my_type==5 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_191.vcd");
  if(my_type==5 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_192.vcd");
  if(my_type==5 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_193.vcd");
  if(my_type==5 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_194.vcd");
  if(my_type==5 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_195.vcd");
  if(my_type==5 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_196.vcd");
  if(my_type==5 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_197.vcd");
  if(my_type==5 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_198.vcd");
  if(my_type==5 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_199.vcd");
  if(my_type==5 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_200.vcd");
  if(my_type==5 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_201.vcd");
  if(my_type==5 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_202.vcd");
  if(my_type==5 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_203.vcd");
  if(my_type==5 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_204.vcd");
  if(my_type==5 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_205.vcd");
  if(my_type==5 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_206.vcd");
  if(my_type==5 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_207.vcd");
  if(my_type==5 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_208.vcd");
  if(my_type==5 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_209.vcd");
  if(my_type==5 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_210.vcd");
  if(my_type==5 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_211.vcd");
  if(my_type==5 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_212.vcd");
  if(my_type==5 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_213.vcd");
  if(my_type==5 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_214.vcd");
  if(my_type==5 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_215.vcd");
  if(my_type==5 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_216.vcd");
  if(my_type==5 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_217.vcd");
  if(my_type==5 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_218.vcd");
  if(my_type==5 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_219.vcd");
  if(my_type==5 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_220.vcd");
  if(my_type==5 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_221.vcd");
  if(my_type==5 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_222.vcd");
  if(my_type==5 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_223.vcd");
  if(my_type==5 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_224.vcd");
  if(my_type==5 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_225.vcd");
  if(my_type==5 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_226.vcd");
  if(my_type==5 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_227.vcd");
  if(my_type==5 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_228.vcd");
  if(my_type==5 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_229.vcd");
  if(my_type==5 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_230.vcd");
  if(my_type==5 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_231.vcd");
  if(my_type==5 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_232.vcd");
  if(my_type==5 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_233.vcd");
  if(my_type==5 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_234.vcd");
  if(my_type==5 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_235.vcd");
  if(my_type==5 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_236.vcd");
  if(my_type==5 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_237.vcd");
  if(my_type==5 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_238.vcd");
  if(my_type==5 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_239.vcd");
  if(my_type==5 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_240.vcd");
  if(my_type==5 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_241.vcd");
  if(my_type==5 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_242.vcd");
  if(my_type==5 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_243.vcd");
  if(my_type==5 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_244.vcd");
  if(my_type==5 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_245.vcd");
  if(my_type==5 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_246.vcd");
  if(my_type==5 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_247.vcd");
  if(my_type==5 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_248.vcd");
  if(my_type==5 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_249.vcd");
  if(my_type==5 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_250.vcd");
  if(my_type==5 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_251.vcd");
  if(my_type==5 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_252.vcd");
  if(my_type==5 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_253.vcd");
  if(my_type==5 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_254.vcd");
  if(my_type==5 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_255.vcd");
  if(my_type==5 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_256.vcd");
  if(my_type==5 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_257.vcd");
  if(my_type==5 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_258.vcd");
  if(my_type==5 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_259.vcd");
  if(my_type==5 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_260.vcd");
  if(my_type==5 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_261.vcd");
  if(my_type==5 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_262.vcd");
  if(my_type==5 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_263.vcd");
  if(my_type==5 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_264.vcd");
  if(my_type==5 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_265.vcd");
  if(my_type==5 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_266.vcd");
  if(my_type==5 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_267.vcd");
  if(my_type==5 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_268.vcd");
  if(my_type==5 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_269.vcd");
  if(my_type==5 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_270.vcd");
  if(my_type==5 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_271.vcd");
  if(my_type==5 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_272.vcd");
  if(my_type==5 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_273.vcd");
  if(my_type==5 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_274.vcd");
  if(my_type==5 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_275.vcd");
  if(my_type==5 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_276.vcd");
  if(my_type==5 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_277.vcd");
  if(my_type==5 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_278.vcd");
  if(my_type==5 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_279.vcd");
  if(my_type==5 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_280.vcd");
  if(my_type==5 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_281.vcd");
  if(my_type==5 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_282.vcd");
  if(my_type==5 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_283.vcd");
  if(my_type==5 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_284.vcd");
  if(my_type==5 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_285.vcd");
  if(my_type==5 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_286.vcd");
  if(my_type==5 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_287.vcd");
  if(my_type==5 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_288.vcd");
  if(my_type==5 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_289.vcd");
  if(my_type==5 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_290.vcd");
  if(my_type==5 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_291.vcd");
  if(my_type==5 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_292.vcd");
  if(my_type==5 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_293.vcd");
  if(my_type==5 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_294.vcd");
  if(my_type==5 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_295.vcd");
  if(my_type==5 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_296.vcd");
  if(my_type==5 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_297.vcd");
  if(my_type==5 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_298.vcd");
  if(my_type==5 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_299.vcd");
  if(my_type==5 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_300.vcd");
  if(my_type==5 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_301.vcd");
  if(my_type==5 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_302.vcd");
  if(my_type==5 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_303.vcd");
  if(my_type==5 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_304.vcd");
  if(my_type==5 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_305.vcd");
  if(my_type==5 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_306.vcd");
  if(my_type==5 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_307.vcd");
  if(my_type==5 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_308.vcd");
  if(my_type==5 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_309.vcd");
  if(my_type==5 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_310.vcd");
  if(my_type==5 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_311.vcd");
  if(my_type==5 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_312.vcd");
  if(my_type==5 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_313.vcd");
  if(my_type==5 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_314.vcd");
  if(my_type==5 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_315.vcd");
  if(my_type==5 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_316.vcd");
  if(my_type==5 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_317.vcd");
  if(my_type==5 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_318.vcd");
  if(my_type==5 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_319.vcd");
  if(my_type==5 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_320.vcd");
  if(my_type==5 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_321.vcd");
  if(my_type==5 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_322.vcd");
  if(my_type==5 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_323.vcd");
  if(my_type==5 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_324.vcd");
  if(my_type==5 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_325.vcd");
  if(my_type==5 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_326.vcd");
  if(my_type==5 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_327.vcd");
  if(my_type==5 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_328.vcd");
  if(my_type==5 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_329.vcd");
  if(my_type==5 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_330.vcd");
  if(my_type==5 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_331.vcd");
  if(my_type==5 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_332.vcd");
  if(my_type==5 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_333.vcd");
  if(my_type==5 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_334.vcd");
  if(my_type==5 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_335.vcd");
  if(my_type==5 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_336.vcd");
  if(my_type==5 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_337.vcd");
  if(my_type==5 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_338.vcd");
  if(my_type==5 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_339.vcd");
  if(my_type==5 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_340.vcd");
  if(my_type==5 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_341.vcd");
  if(my_type==5 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_342.vcd");
  if(my_type==5 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_343.vcd");
  if(my_type==5 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_344.vcd");
  if(my_type==5 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_345.vcd");
  if(my_type==5 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_346.vcd");
  if(my_type==5 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_347.vcd");
  if(my_type==5 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_348.vcd");
  if(my_type==5 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_349.vcd");
  if(my_type==5 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_350.vcd");
  if(my_type==5 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_351.vcd");
  if(my_type==5 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_352.vcd");
  if(my_type==5 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_353.vcd");
  if(my_type==5 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_354.vcd");
  if(my_type==5 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_355.vcd");
  if(my_type==5 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_356.vcd");
  if(my_type==5 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_357.vcd");
  if(my_type==5 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_358.vcd");
  if(my_type==5 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_359.vcd");
  if(my_type==5 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_360.vcd");
  if(my_type==5 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_361.vcd");
  if(my_type==5 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_362.vcd");
  if(my_type==5 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_363.vcd");
  if(my_type==5 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_364.vcd");
  if(my_type==5 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_365.vcd");
  if(my_type==5 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_366.vcd");
  if(my_type==5 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_367.vcd");
  if(my_type==5 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_368.vcd");
  if(my_type==5 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_369.vcd");
  if(my_type==5 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_370.vcd");
  if(my_type==5 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_371.vcd");
  if(my_type==5 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_372.vcd");
  if(my_type==5 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_373.vcd");
  if(my_type==5 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_374.vcd");
  if(my_type==5 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_375.vcd");
  if(my_type==5 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_376.vcd");
  if(my_type==5 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_377.vcd");
  if(my_type==5 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_378.vcd");
  if(my_type==5 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_379.vcd");
  if(my_type==5 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_380.vcd");
  if(my_type==5 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_381.vcd");
  if(my_type==5 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_382.vcd");
  if(my_type==5 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_383.vcd");
  if(my_type==5 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_384.vcd");
  if(my_type==5 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_385.vcd");
  if(my_type==5 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_386.vcd");
  if(my_type==5 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_387.vcd");
  if(my_type==5 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_388.vcd");
  if(my_type==5 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_389.vcd");
  if(my_type==5 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_390.vcd");
  if(my_type==5 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_391.vcd");
  if(my_type==5 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_392.vcd");
  if(my_type==5 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_393.vcd");
  if(my_type==5 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_394.vcd");
  if(my_type==5 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_395.vcd");
  if(my_type==5 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_396.vcd");
  if(my_type==5 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_397.vcd");
  if(my_type==5 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_398.vcd");
  if(my_type==5 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_399.vcd");
  if(my_type==5 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_400.vcd");
  if(my_type==5 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_401.vcd");
  if(my_type==5 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_402.vcd");
  if(my_type==5 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_403.vcd");
  if(my_type==5 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_404.vcd");
  if(my_type==5 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_405.vcd");
  if(my_type==5 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_406.vcd");
  if(my_type==5 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_407.vcd");
  if(my_type==5 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_408.vcd");
  if(my_type==5 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_409.vcd");
  if(my_type==5 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_410.vcd");
  if(my_type==5 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_411.vcd");
  if(my_type==5 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_412.vcd");
  if(my_type==5 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_413.vcd");
  if(my_type==5 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_414.vcd");
  if(my_type==5 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_415.vcd");
  if(my_type==5 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_416.vcd");
  if(my_type==5 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_417.vcd");
  if(my_type==5 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_418.vcd");
  if(my_type==5 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_419.vcd");
  if(my_type==5 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_420.vcd");
  if(my_type==5 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_421.vcd");
  if(my_type==5 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_422.vcd");
  if(my_type==5 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_423.vcd");
  if(my_type==5 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_424.vcd");
  if(my_type==5 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_425.vcd");
  if(my_type==5 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_426.vcd");
  if(my_type==5 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_427.vcd");
  if(my_type==5 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_428.vcd");
  if(my_type==5 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_429.vcd");
  if(my_type==5 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_430.vcd");
  if(my_type==5 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_431.vcd");
  if(my_type==5 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_432.vcd");
  if(my_type==5 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_433.vcd");
  if(my_type==5 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_434.vcd");
  if(my_type==5 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_435.vcd");
  if(my_type==5 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_436.vcd");
  if(my_type==5 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_437.vcd");
  if(my_type==5 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_438.vcd");
  if(my_type==5 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_439.vcd");
  if(my_type==5 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_440.vcd");
  if(my_type==5 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_441.vcd");
  if(my_type==5 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_442.vcd");
  if(my_type==5 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_443.vcd");
  if(my_type==5 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_444.vcd");
  if(my_type==5 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_445.vcd");
  if(my_type==5 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_446.vcd");
  if(my_type==5 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_447.vcd");
  if(my_type==5 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_448.vcd");
  if(my_type==5 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_449.vcd");
  if(my_type==5 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_450.vcd");
  if(my_type==5 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_451.vcd");
  if(my_type==5 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_452.vcd");
  if(my_type==5 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_453.vcd");
  if(my_type==5 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_454.vcd");
  if(my_type==5 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_455.vcd");
  if(my_type==5 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_456.vcd");
  if(my_type==5 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_457.vcd");
  if(my_type==5 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_458.vcd");
  if(my_type==5 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_459.vcd");
  if(my_type==5 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_460.vcd");
  if(my_type==5 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_461.vcd");
  if(my_type==5 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_462.vcd");
  if(my_type==5 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_463.vcd");
  if(my_type==5 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_464.vcd");
  if(my_type==5 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_465.vcd");
  if(my_type==5 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_466.vcd");
  if(my_type==5 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_467.vcd");
  if(my_type==5 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_468.vcd");
  if(my_type==5 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_469.vcd");
  if(my_type==5 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_470.vcd");
  if(my_type==5 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_471.vcd");
  if(my_type==5 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_472.vcd");
  if(my_type==5 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_473.vcd");
  if(my_type==5 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_474.vcd");
  if(my_type==5 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_475.vcd");
  if(my_type==5 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_476.vcd");
  if(my_type==5 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_477.vcd");
  if(my_type==5 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_478.vcd");
  if(my_type==5 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_479.vcd");
  if(my_type==5 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_480.vcd");
  if(my_type==5 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_481.vcd");
  if(my_type==5 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_482.vcd");
  if(my_type==5 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_483.vcd");
  if(my_type==5 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_484.vcd");
  if(my_type==5 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_485.vcd");
  if(my_type==5 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_486.vcd");
  if(my_type==5 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_487.vcd");
  if(my_type==5 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_488.vcd");
  if(my_type==5 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_489.vcd");
  if(my_type==5 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_490.vcd");
  if(my_type==5 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_491.vcd");
  if(my_type==5 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_492.vcd");
  if(my_type==5 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_493.vcd");
  if(my_type==5 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_494.vcd");
  if(my_type==5 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_495.vcd");
  if(my_type==5 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_496.vcd");
  if(my_type==5 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_497.vcd");
  if(my_type==5 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_498.vcd");
  if(my_type==5 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_499.vcd");
  if(my_type==5 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_500.vcd");
  if(my_type==5 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_501.vcd");
  if(my_type==5 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_502.vcd");
  if(my_type==5 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_503.vcd");
  if(my_type==5 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_504.vcd");
  if(my_type==5 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_505.vcd");
  if(my_type==5 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_506.vcd");
  if(my_type==5 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_507.vcd");
  if(my_type==5 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_508.vcd");
  if(my_type==5 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_509.vcd");
  if(my_type==5 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_510.vcd");
  if(my_type==5 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_511.vcd");
  if(my_type==5 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_512.vcd");
  if(my_type==5 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_513.vcd");
  if(my_type==5 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_514.vcd");
  if(my_type==5 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_515.vcd");
  if(my_type==5 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_516.vcd");
  if(my_type==5 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_517.vcd");
  if(my_type==5 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_518.vcd");
  if(my_type==5 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_519.vcd");
  if(my_type==5 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_520.vcd");
  if(my_type==5 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_521.vcd");
  if(my_type==5 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_522.vcd");
  if(my_type==5 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_523.vcd");
  if(my_type==5 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_524.vcd");
  if(my_type==5 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_525.vcd");
  if(my_type==5 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_526.vcd");
  if(my_type==5 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_527.vcd");
  if(my_type==5 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_528.vcd");
  if(my_type==5 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_529.vcd");
  if(my_type==5 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_530.vcd");
  if(my_type==5 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_531.vcd");
  if(my_type==5 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_532.vcd");
  if(my_type==5 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_533.vcd");
  if(my_type==5 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_534.vcd");
  if(my_type==5 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_535.vcd");
  if(my_type==5 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_536.vcd");
  if(my_type==5 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_537.vcd");
  if(my_type==5 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_538.vcd");
  if(my_type==5 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_539.vcd");
  if(my_type==5 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_540.vcd");
  if(my_type==5 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_541.vcd");
  if(my_type==5 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_542.vcd");
  if(my_type==5 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_543.vcd");
  if(my_type==5 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_544.vcd");
  if(my_type==5 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_545.vcd");
  if(my_type==5 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_546.vcd");
  if(my_type==5 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_547.vcd");
  if(my_type==5 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_548.vcd");
  if(my_type==5 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_549.vcd");
  if(my_type==5 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_550.vcd");
  if(my_type==5 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_551.vcd");
  if(my_type==5 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_552.vcd");
  if(my_type==5 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_553.vcd");
  if(my_type==5 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_554.vcd");
  if(my_type==5 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_555.vcd");
  if(my_type==5 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_556.vcd");
  if(my_type==5 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_557.vcd");
  if(my_type==5 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_558.vcd");
  if(my_type==5 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_559.vcd");
  if(my_type==5 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_560.vcd");
  if(my_type==5 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_561.vcd");
  if(my_type==5 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_562.vcd");
  if(my_type==5 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_563.vcd");
  if(my_type==5 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_564.vcd");
  if(my_type==5 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_565.vcd");
  if(my_type==5 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_566.vcd");
  if(my_type==5 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_567.vcd");
  if(my_type==5 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_568.vcd");
  if(my_type==5 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_569.vcd");
  if(my_type==5 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_570.vcd");
  if(my_type==5 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_571.vcd");
  if(my_type==5 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_572.vcd");
  if(my_type==5 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_573.vcd");
  if(my_type==5 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_574.vcd");
  if(my_type==5 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_575.vcd");
  if(my_type==5 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_576.vcd");
  if(my_type==5 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_577.vcd");
  if(my_type==5 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_578.vcd");
  if(my_type==5 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_579.vcd");
  if(my_type==5 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_580.vcd");
  if(my_type==5 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_581.vcd");
  if(my_type==5 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_582.vcd");
  if(my_type==5 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_583.vcd");
  if(my_type==5 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_584.vcd");
  if(my_type==5 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_585.vcd");
  if(my_type==5 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_586.vcd");
  if(my_type==5 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_587.vcd");
  if(my_type==5 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_588.vcd");
  if(my_type==5 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_589.vcd");
  if(my_type==5 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_590.vcd");
  if(my_type==5 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_591.vcd");
  if(my_type==5 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_592.vcd");
  if(my_type==5 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_593.vcd");
  if(my_type==5 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_594.vcd");
  if(my_type==5 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_595.vcd");
  if(my_type==5 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_596.vcd");
  if(my_type==5 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_597.vcd");
  if(my_type==5 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_598.vcd");
  if(my_type==5 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_599.vcd");
  if(my_type==5 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_600.vcd");
  if(my_type==5 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_601.vcd");
  if(my_type==5 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_602.vcd");
  if(my_type==5 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_603.vcd");
  if(my_type==5 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_604.vcd");
  if(my_type==5 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_605.vcd");
  if(my_type==5 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_606.vcd");
  if(my_type==5 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_607.vcd");
  if(my_type==5 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_608.vcd");
  if(my_type==5 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_609.vcd");
  if(my_type==5 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_610.vcd");
  if(my_type==5 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_611.vcd");
  if(my_type==5 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_612.vcd");
  if(my_type==5 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_613.vcd");
  if(my_type==5 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_614.vcd");
  if(my_type==5 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_615.vcd");
  if(my_type==5 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_616.vcd");
  if(my_type==5 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_617.vcd");
  if(my_type==5 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_618.vcd");
  if(my_type==5 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_619.vcd");
  if(my_type==5 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_620.vcd");
  if(my_type==5 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_621.vcd");
  if(my_type==5 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_622.vcd");
  if(my_type==5 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_623.vcd");
  if(my_type==5 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_624.vcd");
  if(my_type==5 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_625.vcd");
  if(my_type==5 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_626.vcd");
  if(my_type==5 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_627.vcd");
  if(my_type==5 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_628.vcd");
  if(my_type==5 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_629.vcd");
  if(my_type==5 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_630.vcd");
  if(my_type==5 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_631.vcd");
  if(my_type==5 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_632.vcd");
  if(my_type==5 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_633.vcd");
  if(my_type==5 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_634.vcd");
  if(my_type==5 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_635.vcd");
  if(my_type==5 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_636.vcd");
  if(my_type==5 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_637.vcd");
  if(my_type==5 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_638.vcd");
  if(my_type==5 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_639.vcd");
  if(my_type==5 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_640.vcd");
  if(my_type==5 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_641.vcd");
  if(my_type==5 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_642.vcd");
  if(my_type==5 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_643.vcd");
  if(my_type==5 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_644.vcd");
  if(my_type==5 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_645.vcd");
  if(my_type==5 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_646.vcd");
  if(my_type==5 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_647.vcd");
  if(my_type==5 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_648.vcd");
  if(my_type==5 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_649.vcd");
  if(my_type==5 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_650.vcd");
  if(my_type==5 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_651.vcd");
  if(my_type==5 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_652.vcd");
  if(my_type==5 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_653.vcd");
  if(my_type==5 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_654.vcd");
  if(my_type==5 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_655.vcd");
  if(my_type==5 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_656.vcd");
  if(my_type==5 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_657.vcd");
  if(my_type==5 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_658.vcd");
  if(my_type==5 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_659.vcd");
  if(my_type==5 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_660.vcd");
  if(my_type==5 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_661.vcd");
  if(my_type==5 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_662.vcd");
  if(my_type==5 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_663.vcd");
  if(my_type==5 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_664.vcd");
  if(my_type==5 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_665.vcd");
  if(my_type==5 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_666.vcd");
  if(my_type==5 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_667.vcd");
  if(my_type==5 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_668.vcd");
  if(my_type==5 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_669.vcd");
  if(my_type==5 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_670.vcd");
  if(my_type==5 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_671.vcd");
  if(my_type==5 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_672.vcd");
  if(my_type==5 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_673.vcd");
  if(my_type==5 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_674.vcd");
  if(my_type==5 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_675.vcd");
  if(my_type==5 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_676.vcd");
  if(my_type==5 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_677.vcd");
  if(my_type==5 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_678.vcd");
  if(my_type==5 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_679.vcd");
  if(my_type==5 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_680.vcd");
  if(my_type==5 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_681.vcd");
  if(my_type==5 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_682.vcd");
  if(my_type==5 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_683.vcd");
  if(my_type==5 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_684.vcd");
  if(my_type==5 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_685.vcd");
  if(my_type==5 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_686.vcd");
  if(my_type==5 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_687.vcd");
  if(my_type==5 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_688.vcd");
  if(my_type==5 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_689.vcd");
  if(my_type==5 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_690.vcd");
  if(my_type==5 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_691.vcd");
  if(my_type==5 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_692.vcd");
  if(my_type==5 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_693.vcd");
  if(my_type==5 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_694.vcd");
  if(my_type==5 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_695.vcd");
  if(my_type==5 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_696.vcd");
  if(my_type==5 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_697.vcd");
  if(my_type==5 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_698.vcd");
  if(my_type==5 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_699.vcd");
  if(my_type==5 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_700.vcd");
  if(my_type==5 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_701.vcd");
  if(my_type==5 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_702.vcd");
  if(my_type==5 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_703.vcd");
  if(my_type==5 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_704.vcd");
  if(my_type==5 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_705.vcd");
  if(my_type==5 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_706.vcd");
  if(my_type==5 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_707.vcd");
  if(my_type==5 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_708.vcd");
  if(my_type==5 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_709.vcd");
  if(my_type==5 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_710.vcd");
  if(my_type==5 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_711.vcd");
  if(my_type==5 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_712.vcd");
  if(my_type==5 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_713.vcd");
  if(my_type==5 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_714.vcd");
  if(my_type==5 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_715.vcd");
  if(my_type==5 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_716.vcd");
  if(my_type==5 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_717.vcd");
  if(my_type==5 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_718.vcd");
  if(my_type==5 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_719.vcd");
  if(my_type==5 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_720.vcd");
  if(my_type==5 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_721.vcd");
  if(my_type==5 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_722.vcd");
  if(my_type==5 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_723.vcd");
  if(my_type==5 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_724.vcd");
  if(my_type==5 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_725.vcd");
  if(my_type==5 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_726.vcd");
  if(my_type==5 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_727.vcd");
  if(my_type==5 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_728.vcd");
  if(my_type==5 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_729.vcd");
  if(my_type==5 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_730.vcd");
  if(my_type==5 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_731.vcd");
  if(my_type==5 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_732.vcd");
  if(my_type==5 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_733.vcd");
  if(my_type==5 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_734.vcd");
  if(my_type==5 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_735.vcd");
  if(my_type==5 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_736.vcd");
  if(my_type==5 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_737.vcd");
  if(my_type==5 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_738.vcd");
  if(my_type==5 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_739.vcd");
  if(my_type==5 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_740.vcd");
  if(my_type==5 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_741.vcd");
  if(my_type==5 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_742.vcd");
  if(my_type==5 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_743.vcd");
  if(my_type==5 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_744.vcd");
  if(my_type==5 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_745.vcd");
  if(my_type==5 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_746.vcd");
  if(my_type==5 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_747.vcd");
  if(my_type==5 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_748.vcd");
  if(my_type==5 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_749.vcd");
  if(my_type==5 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_750.vcd");
  if(my_type==5 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_751.vcd");
  if(my_type==5 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_752.vcd");
  if(my_type==5 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_753.vcd");
  if(my_type==5 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_754.vcd");
  if(my_type==5 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_755.vcd");
  if(my_type==5 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_756.vcd");
  if(my_type==5 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_757.vcd");
  if(my_type==5 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_758.vcd");
  if(my_type==5 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_759.vcd");
  if(my_type==5 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_760.vcd");
  if(my_type==5 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_761.vcd");
  if(my_type==5 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_762.vcd");
  if(my_type==5 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_763.vcd");
  if(my_type==5 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_764.vcd");
  if(my_type==5 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_765.vcd");
  if(my_type==5 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_766.vcd");
  if(my_type==5 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_767.vcd");
  if(my_type==5 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_768.vcd");
  if(my_type==5 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_769.vcd");
  if(my_type==5 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_770.vcd");
  if(my_type==5 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_771.vcd");
  if(my_type==5 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_772.vcd");
  if(my_type==5 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_773.vcd");
  if(my_type==5 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_774.vcd");
  if(my_type==5 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_775.vcd");
  if(my_type==5 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_776.vcd");
  if(my_type==5 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_777.vcd");
  if(my_type==5 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_778.vcd");
  if(my_type==5 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_779.vcd");
  if(my_type==5 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_780.vcd");
  if(my_type==5 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_781.vcd");
  if(my_type==5 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_782.vcd");
  if(my_type==5 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_783.vcd");
  if(my_type==5 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_784.vcd");
  if(my_type==5 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_785.vcd");
  if(my_type==5 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_786.vcd");
  if(my_type==5 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_787.vcd");
  if(my_type==5 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_788.vcd");
  if(my_type==5 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_789.vcd");
  if(my_type==5 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_790.vcd");
  if(my_type==5 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_791.vcd");
  if(my_type==5 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_792.vcd");
  if(my_type==5 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_793.vcd");
  if(my_type==5 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_794.vcd");
  if(my_type==5 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_795.vcd");
  if(my_type==5 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_796.vcd");
  if(my_type==5 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_797.vcd");
  if(my_type==5 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_798.vcd");
  if(my_type==5 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_799.vcd");
  if(my_type==5 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_800.vcd");
  if(my_type==5 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_801.vcd");
  if(my_type==5 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_802.vcd");
  if(my_type==5 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_803.vcd");
  if(my_type==5 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_804.vcd");
  if(my_type==5 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_805.vcd");
  if(my_type==5 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_806.vcd");
  if(my_type==5 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_807.vcd");
  if(my_type==5 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_808.vcd");
  if(my_type==5 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_809.vcd");
  if(my_type==5 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_810.vcd");
  if(my_type==5 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_811.vcd");
  if(my_type==5 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_812.vcd");
  if(my_type==5 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_813.vcd");
  if(my_type==5 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_814.vcd");
  if(my_type==5 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_815.vcd");
  if(my_type==5 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_816.vcd");
  if(my_type==5 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_817.vcd");
  if(my_type==5 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_818.vcd");
  if(my_type==5 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_819.vcd");
  if(my_type==5 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_820.vcd");
  if(my_type==5 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_821.vcd");
  if(my_type==5 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_822.vcd");
  if(my_type==5 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_823.vcd");
  if(my_type==5 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_824.vcd");
  if(my_type==5 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_825.vcd");
  if(my_type==5 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_826.vcd");
  if(my_type==5 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_827.vcd");
  if(my_type==5 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_828.vcd");
  if(my_type==5 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_829.vcd");
  if(my_type==5 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_830.vcd");
  if(my_type==5 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_831.vcd");
  if(my_type==5 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_832.vcd");
  if(my_type==5 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_833.vcd");
  if(my_type==5 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_834.vcd");
  if(my_type==5 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_835.vcd");
  if(my_type==5 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_836.vcd");
  if(my_type==5 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_837.vcd");
  if(my_type==5 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_838.vcd");
  if(my_type==5 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_839.vcd");
  if(my_type==5 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_840.vcd");
  if(my_type==5 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_841.vcd");
  if(my_type==5 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_842.vcd");
  if(my_type==5 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_843.vcd");
  if(my_type==5 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_844.vcd");
  if(my_type==5 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_845.vcd");
  if(my_type==5 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_846.vcd");
  if(my_type==5 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_847.vcd");
  if(my_type==5 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_848.vcd");
  if(my_type==5 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_849.vcd");
  if(my_type==5 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_850.vcd");
  if(my_type==5 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_851.vcd");
  if(my_type==5 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_852.vcd");
  if(my_type==5 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_853.vcd");
  if(my_type==5 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_854.vcd");
  if(my_type==5 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_855.vcd");
  if(my_type==5 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_856.vcd");
  if(my_type==5 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_857.vcd");
  if(my_type==5 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_858.vcd");
  if(my_type==5 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_859.vcd");
  if(my_type==5 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_860.vcd");
  if(my_type==5 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_861.vcd");
  if(my_type==5 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_862.vcd");
  if(my_type==5 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_863.vcd");
  if(my_type==5 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_864.vcd");
  if(my_type==5 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_865.vcd");
  if(my_type==5 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_866.vcd");
  if(my_type==5 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_867.vcd");
  if(my_type==5 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_868.vcd");
  if(my_type==5 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_869.vcd");
  if(my_type==5 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_870.vcd");
  if(my_type==5 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_871.vcd");
  if(my_type==5 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_872.vcd");
  if(my_type==5 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_873.vcd");
  if(my_type==5 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_874.vcd");
  if(my_type==5 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_875.vcd");
  if(my_type==5 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_876.vcd");
  if(my_type==5 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_877.vcd");
  if(my_type==5 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_878.vcd");
  if(my_type==5 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_879.vcd");
  if(my_type==5 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_880.vcd");
  if(my_type==5 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_881.vcd");
  if(my_type==5 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_882.vcd");
  if(my_type==5 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_883.vcd");
  if(my_type==5 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_884.vcd");
  if(my_type==5 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_885.vcd");
  if(my_type==5 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_886.vcd");
  if(my_type==5 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_887.vcd");
  if(my_type==5 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_888.vcd");
  if(my_type==5 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_889.vcd");
  if(my_type==5 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_890.vcd");
  if(my_type==5 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_891.vcd");
  if(my_type==5 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_892.vcd");
  if(my_type==5 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_893.vcd");
  if(my_type==5 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_894.vcd");
  if(my_type==5 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_895.vcd");
  if(my_type==5 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_896.vcd");
  if(my_type==5 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_897.vcd");
  if(my_type==5 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_898.vcd");
  if(my_type==5 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_899.vcd");
  if(my_type==5 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_900.vcd");
  if(my_type==5 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_901.vcd");
  if(my_type==5 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_902.vcd");
  if(my_type==5 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_903.vcd");
  if(my_type==5 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_904.vcd");
  if(my_type==5 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_905.vcd");
  if(my_type==5 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_906.vcd");
  if(my_type==5 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_907.vcd");
  if(my_type==5 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_908.vcd");
  if(my_type==5 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_909.vcd");
  if(my_type==5 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_910.vcd");
  if(my_type==5 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_911.vcd");
  if(my_type==5 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_912.vcd");
  if(my_type==5 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_913.vcd");
  if(my_type==5 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_914.vcd");
  if(my_type==5 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_915.vcd");
  if(my_type==5 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_916.vcd");
  if(my_type==5 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_917.vcd");
  if(my_type==5 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_918.vcd");
  if(my_type==5 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_919.vcd");
  if(my_type==5 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_920.vcd");
  if(my_type==5 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_921.vcd");
  if(my_type==5 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_922.vcd");
  if(my_type==5 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_923.vcd");
  if(my_type==5 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_924.vcd");
  if(my_type==5 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_925.vcd");
  if(my_type==5 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_926.vcd");
  if(my_type==5 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_927.vcd");
  if(my_type==5 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_928.vcd");
  if(my_type==5 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_929.vcd");
  if(my_type==5 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_930.vcd");
  if(my_type==5 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_931.vcd");
  if(my_type==5 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_932.vcd");
  if(my_type==5 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_933.vcd");
  if(my_type==5 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_934.vcd");
  if(my_type==5 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_935.vcd");
  if(my_type==5 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_936.vcd");
  if(my_type==5 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_937.vcd");
  if(my_type==5 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_938.vcd");
  if(my_type==5 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_939.vcd");
  if(my_type==5 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_940.vcd");
  if(my_type==5 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_941.vcd");
  if(my_type==5 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_942.vcd");
  if(my_type==5 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_943.vcd");
  if(my_type==5 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_944.vcd");
  if(my_type==5 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_945.vcd");
  if(my_type==5 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_946.vcd");
  if(my_type==5 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_947.vcd");
  if(my_type==5 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_948.vcd");
  if(my_type==5 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_949.vcd");
  if(my_type==5 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_950.vcd");
  if(my_type==5 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_951.vcd");
  if(my_type==5 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_952.vcd");
  if(my_type==5 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_953.vcd");
  if(my_type==5 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_954.vcd");
  if(my_type==5 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_955.vcd");
  if(my_type==5 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_956.vcd");
  if(my_type==5 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_957.vcd");
  if(my_type==5 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_958.vcd");
  if(my_type==5 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_959.vcd");
  if(my_type==5 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_960.vcd");
  if(my_type==5 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_961.vcd");
  if(my_type==5 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_962.vcd");
  if(my_type==5 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_963.vcd");
  if(my_type==5 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_964.vcd");
  if(my_type==5 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_965.vcd");
  if(my_type==5 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_966.vcd");
  if(my_type==5 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_967.vcd");
  if(my_type==5 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_968.vcd");
  if(my_type==5 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_969.vcd");
  if(my_type==5 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_970.vcd");
  if(my_type==5 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_971.vcd");
  if(my_type==5 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_972.vcd");
  if(my_type==5 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_973.vcd");
  if(my_type==5 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_974.vcd");
  if(my_type==5 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_975.vcd");
  if(my_type==5 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_976.vcd");
  if(my_type==5 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_977.vcd");
  if(my_type==5 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_978.vcd");
  if(my_type==5 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_979.vcd");
  if(my_type==5 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_980.vcd");
  if(my_type==5 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_981.vcd");
  if(my_type==5 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_982.vcd");
  if(my_type==5 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_983.vcd");
  if(my_type==5 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_984.vcd");
  if(my_type==5 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_985.vcd");
  if(my_type==5 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_986.vcd");
  if(my_type==5 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_987.vcd");
  if(my_type==5 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_988.vcd");
  if(my_type==5 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_989.vcd");
  if(my_type==5 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_990.vcd");
  if(my_type==5 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_991.vcd");
  if(my_type==5 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_992.vcd");
  if(my_type==5 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_993.vcd");
  if(my_type==5 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_994.vcd");
  if(my_type==5 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_995.vcd");
  if(my_type==5 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_996.vcd");
  if(my_type==5 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_997.vcd");
  if(my_type==5 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_998.vcd");
  if(my_type==5 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_5_999.vcd");
  if(my_type==6 && pe_id==0)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_0.vcd");
  if(my_type==6 && pe_id==1)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_1.vcd");
  if(my_type==6 && pe_id==2)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_2.vcd");
  if(my_type==6 && pe_id==3)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_3.vcd");
  if(my_type==6 && pe_id==4)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_4.vcd");
  if(my_type==6 && pe_id==5)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_5.vcd");
  if(my_type==6 && pe_id==6)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_6.vcd");
  if(my_type==6 && pe_id==7)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_7.vcd");
  if(my_type==6 && pe_id==8)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_8.vcd");
  if(my_type==6 && pe_id==9)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_9.vcd");
  if(my_type==6 && pe_id==10)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_10.vcd");
  if(my_type==6 && pe_id==11)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_11.vcd");
  if(my_type==6 && pe_id==12)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_12.vcd");
  if(my_type==6 && pe_id==13)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_13.vcd");
  if(my_type==6 && pe_id==14)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_14.vcd");
  if(my_type==6 && pe_id==15)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_15.vcd");
  if(my_type==6 && pe_id==16)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_16.vcd");
  if(my_type==6 && pe_id==17)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_17.vcd");
  if(my_type==6 && pe_id==18)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_18.vcd");
  if(my_type==6 && pe_id==19)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_19.vcd");
  if(my_type==6 && pe_id==20)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_20.vcd");
  if(my_type==6 && pe_id==21)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_21.vcd");
  if(my_type==6 && pe_id==22)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_22.vcd");
  if(my_type==6 && pe_id==23)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_23.vcd");
  if(my_type==6 && pe_id==24)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_24.vcd");
  if(my_type==6 && pe_id==25)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_25.vcd");
  if(my_type==6 && pe_id==26)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_26.vcd");
  if(my_type==6 && pe_id==27)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_27.vcd");
  if(my_type==6 && pe_id==28)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_28.vcd");
  if(my_type==6 && pe_id==29)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_29.vcd");
  if(my_type==6 && pe_id==30)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_30.vcd");
  if(my_type==6 && pe_id==31)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_31.vcd");
  if(my_type==6 && pe_id==32)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_32.vcd");
  if(my_type==6 && pe_id==33)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_33.vcd");
  if(my_type==6 && pe_id==34)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_34.vcd");
  if(my_type==6 && pe_id==35)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_35.vcd");
  if(my_type==6 && pe_id==36)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_36.vcd");
  if(my_type==6 && pe_id==37)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_37.vcd");
  if(my_type==6 && pe_id==38)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_38.vcd");
  if(my_type==6 && pe_id==39)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_39.vcd");
  if(my_type==6 && pe_id==40)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_40.vcd");
  if(my_type==6 && pe_id==41)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_41.vcd");
  if(my_type==6 && pe_id==42)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_42.vcd");
  if(my_type==6 && pe_id==43)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_43.vcd");
  if(my_type==6 && pe_id==44)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_44.vcd");
  if(my_type==6 && pe_id==45)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_45.vcd");
  if(my_type==6 && pe_id==46)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_46.vcd");
  if(my_type==6 && pe_id==47)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_47.vcd");
  if(my_type==6 && pe_id==48)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_48.vcd");
  if(my_type==6 && pe_id==49)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_49.vcd");
  if(my_type==6 && pe_id==50)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_50.vcd");
  if(my_type==6 && pe_id==51)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_51.vcd");
  if(my_type==6 && pe_id==52)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_52.vcd");
  if(my_type==6 && pe_id==53)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_53.vcd");
  if(my_type==6 && pe_id==54)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_54.vcd");
  if(my_type==6 && pe_id==55)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_55.vcd");
  if(my_type==6 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_56.vcd");
  if(my_type==6 && pe_id==56)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_57.vcd");
  if(my_type==6 && pe_id==58)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_58.vcd");
  if(my_type==6 && pe_id==59)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_59.vcd");
  if(my_type==6 && pe_id==60)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_60.vcd");
  if(my_type==6 && pe_id==61)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_61.vcd");
  if(my_type==6 && pe_id==62)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_62.vcd");
  if(my_type==6 && pe_id==63)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_63.vcd");
  if(my_type==6 && pe_id==64)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_64.vcd");
  if(my_type==6 && pe_id==65)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_65.vcd");
  if(my_type==6 && pe_id==66)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_66.vcd");
  if(my_type==6 && pe_id==67)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_67.vcd");
  if(my_type==6 && pe_id==68)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_68.vcd");
  if(my_type==6 && pe_id==69)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_69.vcd");
  if(my_type==6 && pe_id==70)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_70.vcd");
  if(my_type==6 && pe_id==71)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_71.vcd");
  if(my_type==6 && pe_id==72)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_72.vcd");
  if(my_type==6 && pe_id==73)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_73.vcd");
  if(my_type==6 && pe_id==74)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_74.vcd");
  if(my_type==6 && pe_id==75)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_75.vcd");
  if(my_type==6 && pe_id==76)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_76.vcd");
  if(my_type==6 && pe_id==77)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_77.vcd");
  if(my_type==6 && pe_id==78)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_78.vcd");
  if(my_type==6 && pe_id==79)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_79.vcd");
  if(my_type==6 && pe_id==80)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_80.vcd");
  if(my_type==6 && pe_id==81)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_81.vcd");
  if(my_type==6 && pe_id==82)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_82.vcd");
  if(my_type==6 && pe_id==83)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_83.vcd");
  if(my_type==6 && pe_id==84)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_84.vcd");
  if(my_type==6 && pe_id==85)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_85.vcd");
  if(my_type==6 && pe_id==86)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_86.vcd");
  if(my_type==6 && pe_id==87)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_87.vcd");
  if(my_type==6 && pe_id==88)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_88.vcd");
  if(my_type==6 && pe_id==89)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_89.vcd");
  if(my_type==6 && pe_id==90)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_90.vcd");
  if(my_type==6 && pe_id==91)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_91.vcd");
  if(my_type==6 && pe_id==92)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_92.vcd");
  if(my_type==6 && pe_id==93)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_93.vcd");
  if(my_type==6 && pe_id==94)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_94.vcd");
  if(my_type==6 && pe_id==95)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_95.vcd");
  if(my_type==6 && pe_id==96)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_96.vcd");
  if(my_type==6 && pe_id==97)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_97.vcd");
  if(my_type==6 && pe_id==98)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_98.vcd");
  if(my_type==6 && pe_id==99)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_99.vcd");
  if(my_type==6 && pe_id==100)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_100.vcd");
  if(my_type==6 && pe_id==101)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_101.vcd");
  if(my_type==6 && pe_id==102)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_102.vcd");
  if(my_type==6 && pe_id==103)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_103.vcd");
  if(my_type==6 && pe_id==104)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_104.vcd");
  if(my_type==6 && pe_id==105)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_105.vcd");
  if(my_type==6 && pe_id==106)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_106.vcd");
  if(my_type==6 && pe_id==107)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_107.vcd");
  if(my_type==6 && pe_id==108)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_108.vcd");
  if(my_type==6 && pe_id==109)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_109.vcd");
  if(my_type==6 && pe_id==110)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_110.vcd");
  if(my_type==6 && pe_id==111)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_111.vcd");
  if(my_type==6 && pe_id==112)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_112.vcd");
  if(my_type==6 && pe_id==113)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_113.vcd");
  if(my_type==6 && pe_id==114)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_114.vcd");
  if(my_type==6 && pe_id==115)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_115.vcd");
  if(my_type==6 && pe_id==116)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_116.vcd");
  if(my_type==6 && pe_id==117)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_117.vcd");
  if(my_type==6 && pe_id==118)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_118.vcd");
  if(my_type==6 && pe_id==119)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_119.vcd");
  if(my_type==6 && pe_id==120)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_120.vcd");
  if(my_type==6 && pe_id==121)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_121.vcd");
  if(my_type==6 && pe_id==122)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_122.vcd");
  if(my_type==6 && pe_id==123)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_123.vcd");
  if(my_type==6 && pe_id==124)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_124.vcd");
  if(my_type==6 && pe_id==125)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_125.vcd");
  if(my_type==6 && pe_id==126)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_126.vcd");
  if(my_type==6 && pe_id==127)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_127.vcd");
  if(my_type==6 && pe_id==128)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_128.vcd");
  if(my_type==6 && pe_id==129)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_129.vcd");
  if(my_type==6 && pe_id==130)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_130.vcd");
  if(my_type==6 && pe_id==131)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_131.vcd");
  if(my_type==6 && pe_id==132)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_132.vcd");
  if(my_type==6 && pe_id==133)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_133.vcd");
  if(my_type==6 && pe_id==134)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_134.vcd");
  if(my_type==6 && pe_id==135)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_135.vcd");
  if(my_type==6 && pe_id==136)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_136.vcd");
  if(my_type==6 && pe_id==137)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_137.vcd");
  if(my_type==6 && pe_id==138)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_138.vcd");
  if(my_type==6 && pe_id==139)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_139.vcd");
  if(my_type==6 && pe_id==140)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_140.vcd");
  if(my_type==6 && pe_id==141)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_141.vcd");
  if(my_type==6 && pe_id==142)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_142.vcd");
  if(my_type==6 && pe_id==143)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_143.vcd");
  if(my_type==6 && pe_id==144)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_144.vcd");
  if(my_type==6 && pe_id==145)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_145.vcd");
  if(my_type==6 && pe_id==146)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_146.vcd");
  if(my_type==6 && pe_id==147)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_147.vcd");
  if(my_type==6 && pe_id==148)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_148.vcd");
  if(my_type==6 && pe_id==149)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_149.vcd");
  if(my_type==6 && pe_id==150)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_150.vcd");
  if(my_type==6 && pe_id==151)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_151.vcd");
  if(my_type==6 && pe_id==152)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_152.vcd");
  if(my_type==6 && pe_id==153)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_153.vcd");
  if(my_type==6 && pe_id==154)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_154.vcd");
  if(my_type==6 && pe_id==155)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_155.vcd");
  if(my_type==6 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_156.vcd");
  if(my_type==6 && pe_id==156)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_157.vcd");
  if(my_type==6 && pe_id==158)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_158.vcd");
  if(my_type==6 && pe_id==159)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_159.vcd");
  if(my_type==6 && pe_id==160)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_160.vcd");
  if(my_type==6 && pe_id==161)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_161.vcd");
  if(my_type==6 && pe_id==162)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_162.vcd");
  if(my_type==6 && pe_id==163)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_163.vcd");
  if(my_type==6 && pe_id==164)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_164.vcd");
  if(my_type==6 && pe_id==165)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_165.vcd");
  if(my_type==6 && pe_id==166)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_166.vcd");
  if(my_type==6 && pe_id==167)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_167.vcd");
  if(my_type==6 && pe_id==168)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_168.vcd");
  if(my_type==6 && pe_id==169)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_169.vcd");
  if(my_type==6 && pe_id==170)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_170.vcd");
  if(my_type==6 && pe_id==171)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_171.vcd");
  if(my_type==6 && pe_id==172)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_172.vcd");
  if(my_type==6 && pe_id==173)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_173.vcd");
  if(my_type==6 && pe_id==174)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_174.vcd");
  if(my_type==6 && pe_id==175)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_175.vcd");
  if(my_type==6 && pe_id==176)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_176.vcd");
  if(my_type==6 && pe_id==177)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_177.vcd");
  if(my_type==6 && pe_id==178)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_178.vcd");
  if(my_type==6 && pe_id==179)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_179.vcd");
  if(my_type==6 && pe_id==180)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_180.vcd");
  if(my_type==6 && pe_id==181)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_181.vcd");
  if(my_type==6 && pe_id==182)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_182.vcd");
  if(my_type==6 && pe_id==183)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_183.vcd");
  if(my_type==6 && pe_id==184)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_184.vcd");
  if(my_type==6 && pe_id==185)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_185.vcd");
  if(my_type==6 && pe_id==186)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_186.vcd");
  if(my_type==6 && pe_id==187)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_187.vcd");
  if(my_type==6 && pe_id==188)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_188.vcd");
  if(my_type==6 && pe_id==189)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_189.vcd");
  if(my_type==6 && pe_id==190)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_190.vcd");
  if(my_type==6 && pe_id==191)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_191.vcd");
  if(my_type==6 && pe_id==192)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_192.vcd");
  if(my_type==6 && pe_id==193)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_193.vcd");
  if(my_type==6 && pe_id==194)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_194.vcd");
  if(my_type==6 && pe_id==195)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_195.vcd");
  if(my_type==6 && pe_id==196)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_196.vcd");
  if(my_type==6 && pe_id==197)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_197.vcd");
  if(my_type==6 && pe_id==198)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_198.vcd");
  if(my_type==6 && pe_id==199)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_199.vcd");
  if(my_type==6 && pe_id==200)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_200.vcd");
  if(my_type==6 && pe_id==201)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_201.vcd");
  if(my_type==6 && pe_id==202)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_202.vcd");
  if(my_type==6 && pe_id==203)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_203.vcd");
  if(my_type==6 && pe_id==204)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_204.vcd");
  if(my_type==6 && pe_id==205)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_205.vcd");
  if(my_type==6 && pe_id==206)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_206.vcd");
  if(my_type==6 && pe_id==207)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_207.vcd");
  if(my_type==6 && pe_id==208)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_208.vcd");
  if(my_type==6 && pe_id==209)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_209.vcd");
  if(my_type==6 && pe_id==210)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_210.vcd");
  if(my_type==6 && pe_id==211)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_211.vcd");
  if(my_type==6 && pe_id==212)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_212.vcd");
  if(my_type==6 && pe_id==213)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_213.vcd");
  if(my_type==6 && pe_id==214)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_214.vcd");
  if(my_type==6 && pe_id==215)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_215.vcd");
  if(my_type==6 && pe_id==216)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_216.vcd");
  if(my_type==6 && pe_id==217)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_217.vcd");
  if(my_type==6 && pe_id==218)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_218.vcd");
  if(my_type==6 && pe_id==219)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_219.vcd");
  if(my_type==6 && pe_id==220)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_220.vcd");
  if(my_type==6 && pe_id==221)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_221.vcd");
  if(my_type==6 && pe_id==222)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_222.vcd");
  if(my_type==6 && pe_id==223)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_223.vcd");
  if(my_type==6 && pe_id==224)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_224.vcd");
  if(my_type==6 && pe_id==225)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_225.vcd");
  if(my_type==6 && pe_id==226)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_226.vcd");
  if(my_type==6 && pe_id==227)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_227.vcd");
  if(my_type==6 && pe_id==228)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_228.vcd");
  if(my_type==6 && pe_id==229)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_229.vcd");
  if(my_type==6 && pe_id==230)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_230.vcd");
  if(my_type==6 && pe_id==231)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_231.vcd");
  if(my_type==6 && pe_id==232)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_232.vcd");
  if(my_type==6 && pe_id==233)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_233.vcd");
  if(my_type==6 && pe_id==234)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_234.vcd");
  if(my_type==6 && pe_id==235)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_235.vcd");
  if(my_type==6 && pe_id==236)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_236.vcd");
  if(my_type==6 && pe_id==237)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_237.vcd");
  if(my_type==6 && pe_id==238)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_238.vcd");
  if(my_type==6 && pe_id==239)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_239.vcd");
  if(my_type==6 && pe_id==240)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_240.vcd");
  if(my_type==6 && pe_id==241)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_241.vcd");
  if(my_type==6 && pe_id==242)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_242.vcd");
  if(my_type==6 && pe_id==243)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_243.vcd");
  if(my_type==6 && pe_id==244)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_244.vcd");
  if(my_type==6 && pe_id==245)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_245.vcd");
  if(my_type==6 && pe_id==246)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_246.vcd");
  if(my_type==6 && pe_id==247)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_247.vcd");
  if(my_type==6 && pe_id==248)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_248.vcd");
  if(my_type==6 && pe_id==249)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_249.vcd");
  if(my_type==6 && pe_id==250)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_250.vcd");
  if(my_type==6 && pe_id==251)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_251.vcd");
  if(my_type==6 && pe_id==252)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_252.vcd");
  if(my_type==6 && pe_id==253)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_253.vcd");
  if(my_type==6 && pe_id==254)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_254.vcd");
  if(my_type==6 && pe_id==255)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_255.vcd");
  if(my_type==6 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_256.vcd");
  if(my_type==6 && pe_id==256)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_257.vcd");
  if(my_type==6 && pe_id==258)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_258.vcd");
  if(my_type==6 && pe_id==259)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_259.vcd");
  if(my_type==6 && pe_id==260)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_260.vcd");
  if(my_type==6 && pe_id==261)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_261.vcd");
  if(my_type==6 && pe_id==262)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_262.vcd");
  if(my_type==6 && pe_id==263)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_263.vcd");
  if(my_type==6 && pe_id==264)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_264.vcd");
  if(my_type==6 && pe_id==265)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_265.vcd");
  if(my_type==6 && pe_id==266)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_266.vcd");
  if(my_type==6 && pe_id==267)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_267.vcd");
  if(my_type==6 && pe_id==268)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_268.vcd");
  if(my_type==6 && pe_id==269)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_269.vcd");
  if(my_type==6 && pe_id==270)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_270.vcd");
  if(my_type==6 && pe_id==271)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_271.vcd");
  if(my_type==6 && pe_id==272)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_272.vcd");
  if(my_type==6 && pe_id==273)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_273.vcd");
  if(my_type==6 && pe_id==274)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_274.vcd");
  if(my_type==6 && pe_id==275)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_275.vcd");
  if(my_type==6 && pe_id==276)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_276.vcd");
  if(my_type==6 && pe_id==277)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_277.vcd");
  if(my_type==6 && pe_id==278)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_278.vcd");
  if(my_type==6 && pe_id==279)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_279.vcd");
  if(my_type==6 && pe_id==280)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_280.vcd");
  if(my_type==6 && pe_id==281)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_281.vcd");
  if(my_type==6 && pe_id==282)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_282.vcd");
  if(my_type==6 && pe_id==283)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_283.vcd");
  if(my_type==6 && pe_id==284)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_284.vcd");
  if(my_type==6 && pe_id==285)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_285.vcd");
  if(my_type==6 && pe_id==286)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_286.vcd");
  if(my_type==6 && pe_id==287)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_287.vcd");
  if(my_type==6 && pe_id==288)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_288.vcd");
  if(my_type==6 && pe_id==289)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_289.vcd");
  if(my_type==6 && pe_id==290)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_290.vcd");
  if(my_type==6 && pe_id==291)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_291.vcd");
  if(my_type==6 && pe_id==292)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_292.vcd");
  if(my_type==6 && pe_id==293)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_293.vcd");
  if(my_type==6 && pe_id==294)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_294.vcd");
  if(my_type==6 && pe_id==295)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_295.vcd");
  if(my_type==6 && pe_id==296)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_296.vcd");
  if(my_type==6 && pe_id==297)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_297.vcd");
  if(my_type==6 && pe_id==298)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_298.vcd");
  if(my_type==6 && pe_id==299)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_299.vcd");
  if(my_type==6 && pe_id==300)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_300.vcd");
  if(my_type==6 && pe_id==301)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_301.vcd");
  if(my_type==6 && pe_id==302)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_302.vcd");
  if(my_type==6 && pe_id==303)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_303.vcd");
  if(my_type==6 && pe_id==304)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_304.vcd");
  if(my_type==6 && pe_id==305)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_305.vcd");
  if(my_type==6 && pe_id==306)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_306.vcd");
  if(my_type==6 && pe_id==307)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_307.vcd");
  if(my_type==6 && pe_id==308)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_308.vcd");
  if(my_type==6 && pe_id==309)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_309.vcd");
  if(my_type==6 && pe_id==310)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_310.vcd");
  if(my_type==6 && pe_id==311)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_311.vcd");
  if(my_type==6 && pe_id==312)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_312.vcd");
  if(my_type==6 && pe_id==313)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_313.vcd");
  if(my_type==6 && pe_id==314)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_314.vcd");
  if(my_type==6 && pe_id==315)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_315.vcd");
  if(my_type==6 && pe_id==316)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_316.vcd");
  if(my_type==6 && pe_id==317)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_317.vcd");
  if(my_type==6 && pe_id==318)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_318.vcd");
  if(my_type==6 && pe_id==319)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_319.vcd");
  if(my_type==6 && pe_id==320)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_320.vcd");
  if(my_type==6 && pe_id==321)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_321.vcd");
  if(my_type==6 && pe_id==322)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_322.vcd");
  if(my_type==6 && pe_id==323)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_323.vcd");
  if(my_type==6 && pe_id==324)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_324.vcd");
  if(my_type==6 && pe_id==325)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_325.vcd");
  if(my_type==6 && pe_id==326)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_326.vcd");
  if(my_type==6 && pe_id==327)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_327.vcd");
  if(my_type==6 && pe_id==328)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_328.vcd");
  if(my_type==6 && pe_id==329)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_329.vcd");
  if(my_type==6 && pe_id==330)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_330.vcd");
  if(my_type==6 && pe_id==331)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_331.vcd");
  if(my_type==6 && pe_id==332)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_332.vcd");
  if(my_type==6 && pe_id==333)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_333.vcd");
  if(my_type==6 && pe_id==334)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_334.vcd");
  if(my_type==6 && pe_id==335)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_335.vcd");
  if(my_type==6 && pe_id==336)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_336.vcd");
  if(my_type==6 && pe_id==337)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_337.vcd");
  if(my_type==6 && pe_id==338)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_338.vcd");
  if(my_type==6 && pe_id==339)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_339.vcd");
  if(my_type==6 && pe_id==340)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_340.vcd");
  if(my_type==6 && pe_id==341)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_341.vcd");
  if(my_type==6 && pe_id==342)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_342.vcd");
  if(my_type==6 && pe_id==343)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_343.vcd");
  if(my_type==6 && pe_id==344)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_344.vcd");
  if(my_type==6 && pe_id==345)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_345.vcd");
  if(my_type==6 && pe_id==346)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_346.vcd");
  if(my_type==6 && pe_id==347)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_347.vcd");
  if(my_type==6 && pe_id==348)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_348.vcd");
  if(my_type==6 && pe_id==349)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_349.vcd");
  if(my_type==6 && pe_id==350)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_350.vcd");
  if(my_type==6 && pe_id==351)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_351.vcd");
  if(my_type==6 && pe_id==352)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_352.vcd");
  if(my_type==6 && pe_id==353)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_353.vcd");
  if(my_type==6 && pe_id==354)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_354.vcd");
  if(my_type==6 && pe_id==355)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_355.vcd");
  if(my_type==6 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_356.vcd");
  if(my_type==6 && pe_id==356)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_357.vcd");
  if(my_type==6 && pe_id==358)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_358.vcd");
  if(my_type==6 && pe_id==359)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_359.vcd");
  if(my_type==6 && pe_id==360)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_360.vcd");
  if(my_type==6 && pe_id==361)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_361.vcd");
  if(my_type==6 && pe_id==362)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_362.vcd");
  if(my_type==6 && pe_id==363)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_363.vcd");
  if(my_type==6 && pe_id==364)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_364.vcd");
  if(my_type==6 && pe_id==365)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_365.vcd");
  if(my_type==6 && pe_id==366)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_366.vcd");
  if(my_type==6 && pe_id==367)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_367.vcd");
  if(my_type==6 && pe_id==368)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_368.vcd");
  if(my_type==6 && pe_id==369)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_369.vcd");
  if(my_type==6 && pe_id==370)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_370.vcd");
  if(my_type==6 && pe_id==371)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_371.vcd");
  if(my_type==6 && pe_id==372)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_372.vcd");
  if(my_type==6 && pe_id==373)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_373.vcd");
  if(my_type==6 && pe_id==374)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_374.vcd");
  if(my_type==6 && pe_id==375)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_375.vcd");
  if(my_type==6 && pe_id==376)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_376.vcd");
  if(my_type==6 && pe_id==377)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_377.vcd");
  if(my_type==6 && pe_id==378)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_378.vcd");
  if(my_type==6 && pe_id==379)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_379.vcd");
  if(my_type==6 && pe_id==380)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_380.vcd");
  if(my_type==6 && pe_id==381)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_381.vcd");
  if(my_type==6 && pe_id==382)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_382.vcd");
  if(my_type==6 && pe_id==383)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_383.vcd");
  if(my_type==6 && pe_id==384)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_384.vcd");
  if(my_type==6 && pe_id==385)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_385.vcd");
  if(my_type==6 && pe_id==386)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_386.vcd");
  if(my_type==6 && pe_id==387)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_387.vcd");
  if(my_type==6 && pe_id==388)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_388.vcd");
  if(my_type==6 && pe_id==389)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_389.vcd");
  if(my_type==6 && pe_id==390)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_390.vcd");
  if(my_type==6 && pe_id==391)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_391.vcd");
  if(my_type==6 && pe_id==392)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_392.vcd");
  if(my_type==6 && pe_id==393)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_393.vcd");
  if(my_type==6 && pe_id==394)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_394.vcd");
  if(my_type==6 && pe_id==395)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_395.vcd");
  if(my_type==6 && pe_id==396)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_396.vcd");
  if(my_type==6 && pe_id==397)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_397.vcd");
  if(my_type==6 && pe_id==398)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_398.vcd");
  if(my_type==6 && pe_id==399)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_399.vcd");
  if(my_type==6 && pe_id==400)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_400.vcd");
  if(my_type==6 && pe_id==401)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_401.vcd");
  if(my_type==6 && pe_id==402)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_402.vcd");
  if(my_type==6 && pe_id==403)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_403.vcd");
  if(my_type==6 && pe_id==404)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_404.vcd");
  if(my_type==6 && pe_id==405)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_405.vcd");
  if(my_type==6 && pe_id==406)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_406.vcd");
  if(my_type==6 && pe_id==407)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_407.vcd");
  if(my_type==6 && pe_id==408)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_408.vcd");
  if(my_type==6 && pe_id==409)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_409.vcd");
  if(my_type==6 && pe_id==410)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_410.vcd");
  if(my_type==6 && pe_id==411)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_411.vcd");
  if(my_type==6 && pe_id==412)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_412.vcd");
  if(my_type==6 && pe_id==413)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_413.vcd");
  if(my_type==6 && pe_id==414)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_414.vcd");
  if(my_type==6 && pe_id==415)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_415.vcd");
  if(my_type==6 && pe_id==416)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_416.vcd");
  if(my_type==6 && pe_id==417)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_417.vcd");
  if(my_type==6 && pe_id==418)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_418.vcd");
  if(my_type==6 && pe_id==419)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_419.vcd");
  if(my_type==6 && pe_id==420)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_420.vcd");
  if(my_type==6 && pe_id==421)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_421.vcd");
  if(my_type==6 && pe_id==422)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_422.vcd");
  if(my_type==6 && pe_id==423)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_423.vcd");
  if(my_type==6 && pe_id==424)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_424.vcd");
  if(my_type==6 && pe_id==425)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_425.vcd");
  if(my_type==6 && pe_id==426)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_426.vcd");
  if(my_type==6 && pe_id==427)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_427.vcd");
  if(my_type==6 && pe_id==428)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_428.vcd");
  if(my_type==6 && pe_id==429)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_429.vcd");
  if(my_type==6 && pe_id==430)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_430.vcd");
  if(my_type==6 && pe_id==431)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_431.vcd");
  if(my_type==6 && pe_id==432)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_432.vcd");
  if(my_type==6 && pe_id==433)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_433.vcd");
  if(my_type==6 && pe_id==434)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_434.vcd");
  if(my_type==6 && pe_id==435)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_435.vcd");
  if(my_type==6 && pe_id==436)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_436.vcd");
  if(my_type==6 && pe_id==437)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_437.vcd");
  if(my_type==6 && pe_id==438)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_438.vcd");
  if(my_type==6 && pe_id==439)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_439.vcd");
  if(my_type==6 && pe_id==440)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_440.vcd");
  if(my_type==6 && pe_id==441)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_441.vcd");
  if(my_type==6 && pe_id==442)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_442.vcd");
  if(my_type==6 && pe_id==443)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_443.vcd");
  if(my_type==6 && pe_id==444)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_444.vcd");
  if(my_type==6 && pe_id==445)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_445.vcd");
  if(my_type==6 && pe_id==446)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_446.vcd");
  if(my_type==6 && pe_id==447)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_447.vcd");
  if(my_type==6 && pe_id==448)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_448.vcd");
  if(my_type==6 && pe_id==449)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_449.vcd");
  if(my_type==6 && pe_id==450)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_450.vcd");
  if(my_type==6 && pe_id==451)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_451.vcd");
  if(my_type==6 && pe_id==452)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_452.vcd");
  if(my_type==6 && pe_id==453)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_453.vcd");
  if(my_type==6 && pe_id==454)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_454.vcd");
  if(my_type==6 && pe_id==455)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_455.vcd");
  if(my_type==6 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_456.vcd");
  if(my_type==6 && pe_id==456)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_457.vcd");
  if(my_type==6 && pe_id==458)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_458.vcd");
  if(my_type==6 && pe_id==459)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_459.vcd");
  if(my_type==6 && pe_id==460)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_460.vcd");
  if(my_type==6 && pe_id==461)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_461.vcd");
  if(my_type==6 && pe_id==462)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_462.vcd");
  if(my_type==6 && pe_id==463)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_463.vcd");
  if(my_type==6 && pe_id==464)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_464.vcd");
  if(my_type==6 && pe_id==465)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_465.vcd");
  if(my_type==6 && pe_id==466)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_466.vcd");
  if(my_type==6 && pe_id==467)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_467.vcd");
  if(my_type==6 && pe_id==468)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_468.vcd");
  if(my_type==6 && pe_id==469)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_469.vcd");
  if(my_type==6 && pe_id==470)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_470.vcd");
  if(my_type==6 && pe_id==471)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_471.vcd");
  if(my_type==6 && pe_id==472)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_472.vcd");
  if(my_type==6 && pe_id==473)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_473.vcd");
  if(my_type==6 && pe_id==474)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_474.vcd");
  if(my_type==6 && pe_id==475)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_475.vcd");
  if(my_type==6 && pe_id==476)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_476.vcd");
  if(my_type==6 && pe_id==477)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_477.vcd");
  if(my_type==6 && pe_id==478)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_478.vcd");
  if(my_type==6 && pe_id==479)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_479.vcd");
  if(my_type==6 && pe_id==480)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_480.vcd");
  if(my_type==6 && pe_id==481)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_481.vcd");
  if(my_type==6 && pe_id==482)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_482.vcd");
  if(my_type==6 && pe_id==483)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_483.vcd");
  if(my_type==6 && pe_id==484)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_484.vcd");
  if(my_type==6 && pe_id==485)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_485.vcd");
  if(my_type==6 && pe_id==486)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_486.vcd");
  if(my_type==6 && pe_id==487)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_487.vcd");
  if(my_type==6 && pe_id==488)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_488.vcd");
  if(my_type==6 && pe_id==489)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_489.vcd");
  if(my_type==6 && pe_id==490)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_490.vcd");
  if(my_type==6 && pe_id==491)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_491.vcd");
  if(my_type==6 && pe_id==492)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_492.vcd");
  if(my_type==6 && pe_id==493)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_493.vcd");
  if(my_type==6 && pe_id==494)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_494.vcd");
  if(my_type==6 && pe_id==495)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_495.vcd");
  if(my_type==6 && pe_id==496)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_496.vcd");
  if(my_type==6 && pe_id==497)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_497.vcd");
  if(my_type==6 && pe_id==498)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_498.vcd");
  if(my_type==6 && pe_id==499)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_499.vcd");
  if(my_type==6 && pe_id==500)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_500.vcd");
  if(my_type==6 && pe_id==501)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_501.vcd");
  if(my_type==6 && pe_id==502)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_502.vcd");
  if(my_type==6 && pe_id==503)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_503.vcd");
  if(my_type==6 && pe_id==504)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_504.vcd");
  if(my_type==6 && pe_id==505)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_505.vcd");
  if(my_type==6 && pe_id==506)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_506.vcd");
  if(my_type==6 && pe_id==507)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_507.vcd");
  if(my_type==6 && pe_id==508)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_508.vcd");
  if(my_type==6 && pe_id==509)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_509.vcd");
  if(my_type==6 && pe_id==510)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_510.vcd");
  if(my_type==6 && pe_id==511)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_511.vcd");
  if(my_type==6 && pe_id==512)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_512.vcd");
  if(my_type==6 && pe_id==513)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_513.vcd");
  if(my_type==6 && pe_id==514)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_514.vcd");
  if(my_type==6 && pe_id==515)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_515.vcd");
  if(my_type==6 && pe_id==516)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_516.vcd");
  if(my_type==6 && pe_id==517)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_517.vcd");
  if(my_type==6 && pe_id==518)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_518.vcd");
  if(my_type==6 && pe_id==519)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_519.vcd");
  if(my_type==6 && pe_id==520)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_520.vcd");
  if(my_type==6 && pe_id==521)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_521.vcd");
  if(my_type==6 && pe_id==522)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_522.vcd");
  if(my_type==6 && pe_id==523)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_523.vcd");
  if(my_type==6 && pe_id==524)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_524.vcd");
  if(my_type==6 && pe_id==525)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_525.vcd");
  if(my_type==6 && pe_id==526)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_526.vcd");
  if(my_type==6 && pe_id==527)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_527.vcd");
  if(my_type==6 && pe_id==528)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_528.vcd");
  if(my_type==6 && pe_id==529)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_529.vcd");
  if(my_type==6 && pe_id==530)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_530.vcd");
  if(my_type==6 && pe_id==531)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_531.vcd");
  if(my_type==6 && pe_id==532)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_532.vcd");
  if(my_type==6 && pe_id==533)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_533.vcd");
  if(my_type==6 && pe_id==534)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_534.vcd");
  if(my_type==6 && pe_id==535)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_535.vcd");
  if(my_type==6 && pe_id==536)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_536.vcd");
  if(my_type==6 && pe_id==537)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_537.vcd");
  if(my_type==6 && pe_id==538)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_538.vcd");
  if(my_type==6 && pe_id==539)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_539.vcd");
  if(my_type==6 && pe_id==540)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_540.vcd");
  if(my_type==6 && pe_id==541)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_541.vcd");
  if(my_type==6 && pe_id==542)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_542.vcd");
  if(my_type==6 && pe_id==543)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_543.vcd");
  if(my_type==6 && pe_id==544)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_544.vcd");
  if(my_type==6 && pe_id==545)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_545.vcd");
  if(my_type==6 && pe_id==546)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_546.vcd");
  if(my_type==6 && pe_id==547)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_547.vcd");
  if(my_type==6 && pe_id==548)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_548.vcd");
  if(my_type==6 && pe_id==549)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_549.vcd");
  if(my_type==6 && pe_id==550)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_550.vcd");
  if(my_type==6 && pe_id==551)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_551.vcd");
  if(my_type==6 && pe_id==552)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_552.vcd");
  if(my_type==6 && pe_id==553)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_553.vcd");
  if(my_type==6 && pe_id==554)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_554.vcd");
  if(my_type==6 && pe_id==555)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_555.vcd");
  if(my_type==6 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_556.vcd");
  if(my_type==6 && pe_id==556)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_557.vcd");
  if(my_type==6 && pe_id==558)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_558.vcd");
  if(my_type==6 && pe_id==559)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_559.vcd");
  if(my_type==6 && pe_id==560)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_560.vcd");
  if(my_type==6 && pe_id==561)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_561.vcd");
  if(my_type==6 && pe_id==562)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_562.vcd");
  if(my_type==6 && pe_id==563)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_563.vcd");
  if(my_type==6 && pe_id==564)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_564.vcd");
  if(my_type==6 && pe_id==565)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_565.vcd");
  if(my_type==6 && pe_id==566)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_566.vcd");
  if(my_type==6 && pe_id==567)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_567.vcd");
  if(my_type==6 && pe_id==568)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_568.vcd");
  if(my_type==6 && pe_id==569)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_569.vcd");
  if(my_type==6 && pe_id==570)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_570.vcd");
  if(my_type==6 && pe_id==571)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_571.vcd");
  if(my_type==6 && pe_id==572)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_572.vcd");
  if(my_type==6 && pe_id==573)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_573.vcd");
  if(my_type==6 && pe_id==574)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_574.vcd");
  if(my_type==6 && pe_id==575)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_575.vcd");
  if(my_type==6 && pe_id==576)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_576.vcd");
  if(my_type==6 && pe_id==577)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_577.vcd");
  if(my_type==6 && pe_id==578)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_578.vcd");
  if(my_type==6 && pe_id==579)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_579.vcd");
  if(my_type==6 && pe_id==580)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_580.vcd");
  if(my_type==6 && pe_id==581)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_581.vcd");
  if(my_type==6 && pe_id==582)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_582.vcd");
  if(my_type==6 && pe_id==583)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_583.vcd");
  if(my_type==6 && pe_id==584)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_584.vcd");
  if(my_type==6 && pe_id==585)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_585.vcd");
  if(my_type==6 && pe_id==586)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_586.vcd");
  if(my_type==6 && pe_id==587)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_587.vcd");
  if(my_type==6 && pe_id==588)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_588.vcd");
  if(my_type==6 && pe_id==589)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_589.vcd");
  if(my_type==6 && pe_id==590)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_590.vcd");
  if(my_type==6 && pe_id==591)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_591.vcd");
  if(my_type==6 && pe_id==592)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_592.vcd");
  if(my_type==6 && pe_id==593)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_593.vcd");
  if(my_type==6 && pe_id==594)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_594.vcd");
  if(my_type==6 && pe_id==595)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_595.vcd");
  if(my_type==6 && pe_id==596)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_596.vcd");
  if(my_type==6 && pe_id==597)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_597.vcd");
  if(my_type==6 && pe_id==598)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_598.vcd");
  if(my_type==6 && pe_id==599)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_599.vcd");
  if(my_type==6 && pe_id==600)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_600.vcd");
  if(my_type==6 && pe_id==601)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_601.vcd");
  if(my_type==6 && pe_id==602)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_602.vcd");
  if(my_type==6 && pe_id==603)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_603.vcd");
  if(my_type==6 && pe_id==604)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_604.vcd");
  if(my_type==6 && pe_id==605)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_605.vcd");
  if(my_type==6 && pe_id==606)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_606.vcd");
  if(my_type==6 && pe_id==607)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_607.vcd");
  if(my_type==6 && pe_id==608)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_608.vcd");
  if(my_type==6 && pe_id==609)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_609.vcd");
  if(my_type==6 && pe_id==610)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_610.vcd");
  if(my_type==6 && pe_id==611)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_611.vcd");
  if(my_type==6 && pe_id==612)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_612.vcd");
  if(my_type==6 && pe_id==613)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_613.vcd");
  if(my_type==6 && pe_id==614)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_614.vcd");
  if(my_type==6 && pe_id==615)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_615.vcd");
  if(my_type==6 && pe_id==616)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_616.vcd");
  if(my_type==6 && pe_id==617)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_617.vcd");
  if(my_type==6 && pe_id==618)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_618.vcd");
  if(my_type==6 && pe_id==619)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_619.vcd");
  if(my_type==6 && pe_id==620)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_620.vcd");
  if(my_type==6 && pe_id==621)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_621.vcd");
  if(my_type==6 && pe_id==622)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_622.vcd");
  if(my_type==6 && pe_id==623)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_623.vcd");
  if(my_type==6 && pe_id==624)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_624.vcd");
  if(my_type==6 && pe_id==625)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_625.vcd");
  if(my_type==6 && pe_id==626)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_626.vcd");
  if(my_type==6 && pe_id==627)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_627.vcd");
  if(my_type==6 && pe_id==628)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_628.vcd");
  if(my_type==6 && pe_id==629)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_629.vcd");
  if(my_type==6 && pe_id==630)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_630.vcd");
  if(my_type==6 && pe_id==631)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_631.vcd");
  if(my_type==6 && pe_id==632)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_632.vcd");
  if(my_type==6 && pe_id==633)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_633.vcd");
  if(my_type==6 && pe_id==634)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_634.vcd");
  if(my_type==6 && pe_id==635)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_635.vcd");
  if(my_type==6 && pe_id==636)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_636.vcd");
  if(my_type==6 && pe_id==637)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_637.vcd");
  if(my_type==6 && pe_id==638)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_638.vcd");
  if(my_type==6 && pe_id==639)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_639.vcd");
  if(my_type==6 && pe_id==640)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_640.vcd");
  if(my_type==6 && pe_id==641)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_641.vcd");
  if(my_type==6 && pe_id==642)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_642.vcd");
  if(my_type==6 && pe_id==643)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_643.vcd");
  if(my_type==6 && pe_id==644)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_644.vcd");
  if(my_type==6 && pe_id==645)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_645.vcd");
  if(my_type==6 && pe_id==646)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_646.vcd");
  if(my_type==6 && pe_id==647)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_647.vcd");
  if(my_type==6 && pe_id==648)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_648.vcd");
  if(my_type==6 && pe_id==649)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_649.vcd");
  if(my_type==6 && pe_id==650)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_650.vcd");
  if(my_type==6 && pe_id==651)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_651.vcd");
  if(my_type==6 && pe_id==652)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_652.vcd");
  if(my_type==6 && pe_id==653)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_653.vcd");
  if(my_type==6 && pe_id==654)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_654.vcd");
  if(my_type==6 && pe_id==655)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_655.vcd");
  if(my_type==6 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_656.vcd");
  if(my_type==6 && pe_id==656)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_657.vcd");
  if(my_type==6 && pe_id==658)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_658.vcd");
  if(my_type==6 && pe_id==659)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_659.vcd");
  if(my_type==6 && pe_id==660)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_660.vcd");
  if(my_type==6 && pe_id==661)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_661.vcd");
  if(my_type==6 && pe_id==662)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_662.vcd");
  if(my_type==6 && pe_id==663)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_663.vcd");
  if(my_type==6 && pe_id==664)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_664.vcd");
  if(my_type==6 && pe_id==665)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_665.vcd");
  if(my_type==6 && pe_id==666)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_666.vcd");
  if(my_type==6 && pe_id==667)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_667.vcd");
  if(my_type==6 && pe_id==668)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_668.vcd");
  if(my_type==6 && pe_id==669)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_669.vcd");
  if(my_type==6 && pe_id==670)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_670.vcd");
  if(my_type==6 && pe_id==671)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_671.vcd");
  if(my_type==6 && pe_id==672)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_672.vcd");
  if(my_type==6 && pe_id==673)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_673.vcd");
  if(my_type==6 && pe_id==674)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_674.vcd");
  if(my_type==6 && pe_id==675)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_675.vcd");
  if(my_type==6 && pe_id==676)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_676.vcd");
  if(my_type==6 && pe_id==677)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_677.vcd");
  if(my_type==6 && pe_id==678)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_678.vcd");
  if(my_type==6 && pe_id==679)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_679.vcd");
  if(my_type==6 && pe_id==680)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_680.vcd");
  if(my_type==6 && pe_id==681)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_681.vcd");
  if(my_type==6 && pe_id==682)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_682.vcd");
  if(my_type==6 && pe_id==683)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_683.vcd");
  if(my_type==6 && pe_id==684)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_684.vcd");
  if(my_type==6 && pe_id==685)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_685.vcd");
  if(my_type==6 && pe_id==686)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_686.vcd");
  if(my_type==6 && pe_id==687)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_687.vcd");
  if(my_type==6 && pe_id==688)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_688.vcd");
  if(my_type==6 && pe_id==689)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_689.vcd");
  if(my_type==6 && pe_id==690)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_690.vcd");
  if(my_type==6 && pe_id==691)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_691.vcd");
  if(my_type==6 && pe_id==692)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_692.vcd");
  if(my_type==6 && pe_id==693)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_693.vcd");
  if(my_type==6 && pe_id==694)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_694.vcd");
  if(my_type==6 && pe_id==695)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_695.vcd");
  if(my_type==6 && pe_id==696)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_696.vcd");
  if(my_type==6 && pe_id==697)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_697.vcd");
  if(my_type==6 && pe_id==698)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_698.vcd");
  if(my_type==6 && pe_id==699)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_699.vcd");
  if(my_type==6 && pe_id==700)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_700.vcd");
  if(my_type==6 && pe_id==701)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_701.vcd");
  if(my_type==6 && pe_id==702)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_702.vcd");
  if(my_type==6 && pe_id==703)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_703.vcd");
  if(my_type==6 && pe_id==704)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_704.vcd");
  if(my_type==6 && pe_id==705)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_705.vcd");
  if(my_type==6 && pe_id==706)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_706.vcd");
  if(my_type==6 && pe_id==707)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_707.vcd");
  if(my_type==6 && pe_id==708)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_708.vcd");
  if(my_type==6 && pe_id==709)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_709.vcd");
  if(my_type==6 && pe_id==710)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_710.vcd");
  if(my_type==6 && pe_id==711)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_711.vcd");
  if(my_type==6 && pe_id==712)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_712.vcd");
  if(my_type==6 && pe_id==713)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_713.vcd");
  if(my_type==6 && pe_id==714)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_714.vcd");
  if(my_type==6 && pe_id==715)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_715.vcd");
  if(my_type==6 && pe_id==716)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_716.vcd");
  if(my_type==6 && pe_id==717)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_717.vcd");
  if(my_type==6 && pe_id==718)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_718.vcd");
  if(my_type==6 && pe_id==719)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_719.vcd");
  if(my_type==6 && pe_id==720)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_720.vcd");
  if(my_type==6 && pe_id==721)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_721.vcd");
  if(my_type==6 && pe_id==722)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_722.vcd");
  if(my_type==6 && pe_id==723)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_723.vcd");
  if(my_type==6 && pe_id==724)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_724.vcd");
  if(my_type==6 && pe_id==725)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_725.vcd");
  if(my_type==6 && pe_id==726)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_726.vcd");
  if(my_type==6 && pe_id==727)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_727.vcd");
  if(my_type==6 && pe_id==728)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_728.vcd");
  if(my_type==6 && pe_id==729)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_729.vcd");
  if(my_type==6 && pe_id==730)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_730.vcd");
  if(my_type==6 && pe_id==731)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_731.vcd");
  if(my_type==6 && pe_id==732)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_732.vcd");
  if(my_type==6 && pe_id==733)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_733.vcd");
  if(my_type==6 && pe_id==734)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_734.vcd");
  if(my_type==6 && pe_id==735)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_735.vcd");
  if(my_type==6 && pe_id==736)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_736.vcd");
  if(my_type==6 && pe_id==737)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_737.vcd");
  if(my_type==6 && pe_id==738)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_738.vcd");
  if(my_type==6 && pe_id==739)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_739.vcd");
  if(my_type==6 && pe_id==740)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_740.vcd");
  if(my_type==6 && pe_id==741)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_741.vcd");
  if(my_type==6 && pe_id==742)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_742.vcd");
  if(my_type==6 && pe_id==743)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_743.vcd");
  if(my_type==6 && pe_id==744)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_744.vcd");
  if(my_type==6 && pe_id==745)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_745.vcd");
  if(my_type==6 && pe_id==746)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_746.vcd");
  if(my_type==6 && pe_id==747)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_747.vcd");
  if(my_type==6 && pe_id==748)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_748.vcd");
  if(my_type==6 && pe_id==749)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_749.vcd");
  if(my_type==6 && pe_id==750)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_750.vcd");
  if(my_type==6 && pe_id==751)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_751.vcd");
  if(my_type==6 && pe_id==752)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_752.vcd");
  if(my_type==6 && pe_id==753)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_753.vcd");
  if(my_type==6 && pe_id==754)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_754.vcd");
  if(my_type==6 && pe_id==755)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_755.vcd");
  if(my_type==6 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_756.vcd");
  if(my_type==6 && pe_id==756)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_757.vcd");
  if(my_type==6 && pe_id==758)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_758.vcd");
  if(my_type==6 && pe_id==759)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_759.vcd");
  if(my_type==6 && pe_id==760)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_760.vcd");
  if(my_type==6 && pe_id==761)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_761.vcd");
  if(my_type==6 && pe_id==762)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_762.vcd");
  if(my_type==6 && pe_id==763)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_763.vcd");
  if(my_type==6 && pe_id==764)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_764.vcd");
  if(my_type==6 && pe_id==765)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_765.vcd");
  if(my_type==6 && pe_id==766)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_766.vcd");
  if(my_type==6 && pe_id==767)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_767.vcd");
  if(my_type==6 && pe_id==768)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_768.vcd");
  if(my_type==6 && pe_id==769)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_769.vcd");
  if(my_type==6 && pe_id==770)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_770.vcd");
  if(my_type==6 && pe_id==771)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_771.vcd");
  if(my_type==6 && pe_id==772)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_772.vcd");
  if(my_type==6 && pe_id==773)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_773.vcd");
  if(my_type==6 && pe_id==774)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_774.vcd");
  if(my_type==6 && pe_id==775)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_775.vcd");
  if(my_type==6 && pe_id==776)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_776.vcd");
  if(my_type==6 && pe_id==777)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_777.vcd");
  if(my_type==6 && pe_id==778)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_778.vcd");
  if(my_type==6 && pe_id==779)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_779.vcd");
  if(my_type==6 && pe_id==780)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_780.vcd");
  if(my_type==6 && pe_id==781)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_781.vcd");
  if(my_type==6 && pe_id==782)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_782.vcd");
  if(my_type==6 && pe_id==783)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_783.vcd");
  if(my_type==6 && pe_id==784)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_784.vcd");
  if(my_type==6 && pe_id==785)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_785.vcd");
  if(my_type==6 && pe_id==786)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_786.vcd");
  if(my_type==6 && pe_id==787)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_787.vcd");
  if(my_type==6 && pe_id==788)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_788.vcd");
  if(my_type==6 && pe_id==789)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_789.vcd");
  if(my_type==6 && pe_id==790)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_790.vcd");
  if(my_type==6 && pe_id==791)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_791.vcd");
  if(my_type==6 && pe_id==792)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_792.vcd");
  if(my_type==6 && pe_id==793)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_793.vcd");
  if(my_type==6 && pe_id==794)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_794.vcd");
  if(my_type==6 && pe_id==795)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_795.vcd");
  if(my_type==6 && pe_id==796)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_796.vcd");
  if(my_type==6 && pe_id==797)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_797.vcd");
  if(my_type==6 && pe_id==798)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_798.vcd");
  if(my_type==6 && pe_id==799)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_799.vcd");
  if(my_type==6 && pe_id==800)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_800.vcd");
  if(my_type==6 && pe_id==801)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_801.vcd");
  if(my_type==6 && pe_id==802)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_802.vcd");
  if(my_type==6 && pe_id==803)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_803.vcd");
  if(my_type==6 && pe_id==804)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_804.vcd");
  if(my_type==6 && pe_id==805)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_805.vcd");
  if(my_type==6 && pe_id==806)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_806.vcd");
  if(my_type==6 && pe_id==807)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_807.vcd");
  if(my_type==6 && pe_id==808)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_808.vcd");
  if(my_type==6 && pe_id==809)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_809.vcd");
  if(my_type==6 && pe_id==810)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_810.vcd");
  if(my_type==6 && pe_id==811)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_811.vcd");
  if(my_type==6 && pe_id==812)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_812.vcd");
  if(my_type==6 && pe_id==813)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_813.vcd");
  if(my_type==6 && pe_id==814)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_814.vcd");
  if(my_type==6 && pe_id==815)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_815.vcd");
  if(my_type==6 && pe_id==816)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_816.vcd");
  if(my_type==6 && pe_id==817)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_817.vcd");
  if(my_type==6 && pe_id==818)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_818.vcd");
  if(my_type==6 && pe_id==819)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_819.vcd");
  if(my_type==6 && pe_id==820)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_820.vcd");
  if(my_type==6 && pe_id==821)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_821.vcd");
  if(my_type==6 && pe_id==822)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_822.vcd");
  if(my_type==6 && pe_id==823)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_823.vcd");
  if(my_type==6 && pe_id==824)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_824.vcd");
  if(my_type==6 && pe_id==825)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_825.vcd");
  if(my_type==6 && pe_id==826)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_826.vcd");
  if(my_type==6 && pe_id==827)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_827.vcd");
  if(my_type==6 && pe_id==828)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_828.vcd");
  if(my_type==6 && pe_id==829)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_829.vcd");
  if(my_type==6 && pe_id==830)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_830.vcd");
  if(my_type==6 && pe_id==831)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_831.vcd");
  if(my_type==6 && pe_id==832)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_832.vcd");
  if(my_type==6 && pe_id==833)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_833.vcd");
  if(my_type==6 && pe_id==834)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_834.vcd");
  if(my_type==6 && pe_id==835)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_835.vcd");
  if(my_type==6 && pe_id==836)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_836.vcd");
  if(my_type==6 && pe_id==837)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_837.vcd");
  if(my_type==6 && pe_id==838)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_838.vcd");
  if(my_type==6 && pe_id==839)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_839.vcd");
  if(my_type==6 && pe_id==840)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_840.vcd");
  if(my_type==6 && pe_id==841)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_841.vcd");
  if(my_type==6 && pe_id==842)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_842.vcd");
  if(my_type==6 && pe_id==843)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_843.vcd");
  if(my_type==6 && pe_id==844)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_844.vcd");
  if(my_type==6 && pe_id==845)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_845.vcd");
  if(my_type==6 && pe_id==846)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_846.vcd");
  if(my_type==6 && pe_id==847)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_847.vcd");
  if(my_type==6 && pe_id==848)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_848.vcd");
  if(my_type==6 && pe_id==849)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_849.vcd");
  if(my_type==6 && pe_id==850)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_850.vcd");
  if(my_type==6 && pe_id==851)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_851.vcd");
  if(my_type==6 && pe_id==852)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_852.vcd");
  if(my_type==6 && pe_id==853)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_853.vcd");
  if(my_type==6 && pe_id==854)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_854.vcd");
  if(my_type==6 && pe_id==855)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_855.vcd");
  if(my_type==6 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_856.vcd");
  if(my_type==6 && pe_id==856)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_857.vcd");
  if(my_type==6 && pe_id==858)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_858.vcd");
  if(my_type==6 && pe_id==859)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_859.vcd");
  if(my_type==6 && pe_id==860)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_860.vcd");
  if(my_type==6 && pe_id==861)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_861.vcd");
  if(my_type==6 && pe_id==862)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_862.vcd");
  if(my_type==6 && pe_id==863)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_863.vcd");
  if(my_type==6 && pe_id==864)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_864.vcd");
  if(my_type==6 && pe_id==865)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_865.vcd");
  if(my_type==6 && pe_id==866)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_866.vcd");
  if(my_type==6 && pe_id==867)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_867.vcd");
  if(my_type==6 && pe_id==868)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_868.vcd");
  if(my_type==6 && pe_id==869)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_869.vcd");
  if(my_type==6 && pe_id==870)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_870.vcd");
  if(my_type==6 && pe_id==871)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_871.vcd");
  if(my_type==6 && pe_id==872)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_872.vcd");
  if(my_type==6 && pe_id==873)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_873.vcd");
  if(my_type==6 && pe_id==874)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_874.vcd");
  if(my_type==6 && pe_id==875)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_875.vcd");
  if(my_type==6 && pe_id==876)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_876.vcd");
  if(my_type==6 && pe_id==877)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_877.vcd");
  if(my_type==6 && pe_id==878)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_878.vcd");
  if(my_type==6 && pe_id==879)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_879.vcd");
  if(my_type==6 && pe_id==880)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_880.vcd");
  if(my_type==6 && pe_id==881)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_881.vcd");
  if(my_type==6 && pe_id==882)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_882.vcd");
  if(my_type==6 && pe_id==883)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_883.vcd");
  if(my_type==6 && pe_id==884)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_884.vcd");
  if(my_type==6 && pe_id==885)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_885.vcd");
  if(my_type==6 && pe_id==886)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_886.vcd");
  if(my_type==6 && pe_id==887)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_887.vcd");
  if(my_type==6 && pe_id==888)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_888.vcd");
  if(my_type==6 && pe_id==889)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_889.vcd");
  if(my_type==6 && pe_id==890)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_890.vcd");
  if(my_type==6 && pe_id==891)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_891.vcd");
  if(my_type==6 && pe_id==892)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_892.vcd");
  if(my_type==6 && pe_id==893)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_893.vcd");
  if(my_type==6 && pe_id==894)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_894.vcd");
  if(my_type==6 && pe_id==895)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_895.vcd");
  if(my_type==6 && pe_id==896)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_896.vcd");
  if(my_type==6 && pe_id==897)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_897.vcd");
  if(my_type==6 && pe_id==898)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_898.vcd");
  if(my_type==6 && pe_id==899)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_899.vcd");
  if(my_type==6 && pe_id==900)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_900.vcd");
  if(my_type==6 && pe_id==901)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_901.vcd");
  if(my_type==6 && pe_id==902)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_902.vcd");
  if(my_type==6 && pe_id==903)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_903.vcd");
  if(my_type==6 && pe_id==904)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_904.vcd");
  if(my_type==6 && pe_id==905)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_905.vcd");
  if(my_type==6 && pe_id==906)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_906.vcd");
  if(my_type==6 && pe_id==907)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_907.vcd");
  if(my_type==6 && pe_id==908)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_908.vcd");
  if(my_type==6 && pe_id==909)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_909.vcd");
  if(my_type==6 && pe_id==910)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_910.vcd");
  if(my_type==6 && pe_id==911)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_911.vcd");
  if(my_type==6 && pe_id==912)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_912.vcd");
  if(my_type==6 && pe_id==913)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_913.vcd");
  if(my_type==6 && pe_id==914)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_914.vcd");
  if(my_type==6 && pe_id==915)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_915.vcd");
  if(my_type==6 && pe_id==916)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_916.vcd");
  if(my_type==6 && pe_id==917)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_917.vcd");
  if(my_type==6 && pe_id==918)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_918.vcd");
  if(my_type==6 && pe_id==919)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_919.vcd");
  if(my_type==6 && pe_id==920)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_920.vcd");
  if(my_type==6 && pe_id==921)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_921.vcd");
  if(my_type==6 && pe_id==922)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_922.vcd");
  if(my_type==6 && pe_id==923)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_923.vcd");
  if(my_type==6 && pe_id==924)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_924.vcd");
  if(my_type==6 && pe_id==925)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_925.vcd");
  if(my_type==6 && pe_id==926)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_926.vcd");
  if(my_type==6 && pe_id==927)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_927.vcd");
  if(my_type==6 && pe_id==928)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_928.vcd");
  if(my_type==6 && pe_id==929)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_929.vcd");
  if(my_type==6 && pe_id==930)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_930.vcd");
  if(my_type==6 && pe_id==931)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_931.vcd");
  if(my_type==6 && pe_id==932)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_932.vcd");
  if(my_type==6 && pe_id==933)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_933.vcd");
  if(my_type==6 && pe_id==934)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_934.vcd");
  if(my_type==6 && pe_id==935)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_935.vcd");
  if(my_type==6 && pe_id==936)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_936.vcd");
  if(my_type==6 && pe_id==937)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_937.vcd");
  if(my_type==6 && pe_id==938)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_938.vcd");
  if(my_type==6 && pe_id==939)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_939.vcd");
  if(my_type==6 && pe_id==940)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_940.vcd");
  if(my_type==6 && pe_id==941)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_941.vcd");
  if(my_type==6 && pe_id==942)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_942.vcd");
  if(my_type==6 && pe_id==943)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_943.vcd");
  if(my_type==6 && pe_id==944)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_944.vcd");
  if(my_type==6 && pe_id==945)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_945.vcd");
  if(my_type==6 && pe_id==946)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_946.vcd");
  if(my_type==6 && pe_id==947)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_947.vcd");
  if(my_type==6 && pe_id==948)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_948.vcd");
  if(my_type==6 && pe_id==949)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_949.vcd");
  if(my_type==6 && pe_id==950)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_950.vcd");
  if(my_type==6 && pe_id==951)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_951.vcd");
  if(my_type==6 && pe_id==952)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_952.vcd");
  if(my_type==6 && pe_id==953)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_953.vcd");
  if(my_type==6 && pe_id==954)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_954.vcd");
  if(my_type==6 && pe_id==955)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_955.vcd");
  if(my_type==6 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_956.vcd");
  if(my_type==6 && pe_id==956)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_957.vcd");
  if(my_type==6 && pe_id==958)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_958.vcd");
  if(my_type==6 && pe_id==959)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_959.vcd");
  if(my_type==6 && pe_id==960)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_960.vcd");
  if(my_type==6 && pe_id==961)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_961.vcd");
  if(my_type==6 && pe_id==962)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_962.vcd");
  if(my_type==6 && pe_id==963)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_963.vcd");
  if(my_type==6 && pe_id==964)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_964.vcd");
  if(my_type==6 && pe_id==965)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_965.vcd");
  if(my_type==6 && pe_id==966)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_966.vcd");
  if(my_type==6 && pe_id==967)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_967.vcd");
  if(my_type==6 && pe_id==968)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_968.vcd");
  if(my_type==6 && pe_id==969)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_969.vcd");
  if(my_type==6 && pe_id==970)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_970.vcd");
  if(my_type==6 && pe_id==971)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_971.vcd");
  if(my_type==6 && pe_id==972)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_972.vcd");
  if(my_type==6 && pe_id==973)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_973.vcd");
  if(my_type==6 && pe_id==974)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_974.vcd");
  if(my_type==6 && pe_id==975)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_975.vcd");
  if(my_type==6 && pe_id==976)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_976.vcd");
  if(my_type==6 && pe_id==977)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_977.vcd");
  if(my_type==6 && pe_id==978)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_978.vcd");
  if(my_type==6 && pe_id==979)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_979.vcd");
  if(my_type==6 && pe_id==980)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_980.vcd");
  if(my_type==6 && pe_id==981)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_981.vcd");
  if(my_type==6 && pe_id==982)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_982.vcd");
  if(my_type==6 && pe_id==983)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_983.vcd");
  if(my_type==6 && pe_id==984)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_984.vcd");
  if(my_type==6 && pe_id==985)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_985.vcd");
  if(my_type==6 && pe_id==986)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_986.vcd");
  if(my_type==6 && pe_id==987)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_987.vcd");
  if(my_type==6 && pe_id==988)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_988.vcd");
  if(my_type==6 && pe_id==989)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_989.vcd");
  if(my_type==6 && pe_id==990)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_990.vcd");
  if(my_type==6 && pe_id==991)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_991.vcd");
  if(my_type==6 && pe_id==992)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_992.vcd");
  if(my_type==6 && pe_id==993)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_993.vcd");
  if(my_type==6 && pe_id==994)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_994.vcd");
  if(my_type==6 && pe_id==995)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_995.vcd");
  if(my_type==6 && pe_id==996)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_996.vcd");
  if(my_type==6 && pe_id==997)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_997.vcd");
  if(my_type==6 && pe_id==998)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_998.vcd");
  if(my_type==6 && pe_id==999)$fdumpvars(2,sv_router.router_cortex,"./dump_files/router_6_999.vcd");
  if(my_type>7) $display("Max router's types is 6(0-6)");
  if(pe_id>1000)$display("Max number of routers is 1000(0-999)"); 
 end

endmodule