module router_type_0_netlist;

endmodule