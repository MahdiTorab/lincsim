module router_type_7_netlist;

endmodule