module router_type_1_netlist;

endmodule