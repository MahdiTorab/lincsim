module router_type_5_netlist;

endmodule