module fork_module_netlist;
endmodule