module router_type_4_netlist;

endmodule